VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sram_39_4096
  CLASS BLOCK ;
  FOREIGN sram_39_4096 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1050.000 BY 1600.000 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.040 371.460 97.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.040 371.460 127.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 156.040 371.460 157.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 186.040 371.460 187.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 216.040 371.460 217.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.040 371.460 247.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 276.040 371.460 277.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 306.040 371.460 307.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 336.040 371.460 337.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 366.040 371.460 367.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.040 371.460 397.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 426.040 371.460 427.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 456.040 371.460 457.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 486.040 371.460 487.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 516.040 371.460 517.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.040 371.460 547.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 576.040 371.460 577.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 606.040 371.460 607.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.040 371.460 637.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 666.040 371.460 667.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.040 371.460 697.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 726.040 371.460 727.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 756.040 371.460 757.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.040 371.460 787.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.040 371.460 817.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.040 371.460 847.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 876.040 371.460 877.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 906.040 371.460 907.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 936.040 371.460 937.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 966.040 371.460 967.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.040 371.460 997.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1026.040 371.460 1027.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.040 1168.960 97.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.040 1168.960 127.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 156.040 1168.960 157.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 186.040 1168.960 187.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 216.040 1168.960 217.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.040 1168.960 247.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 276.040 1168.960 277.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 306.040 1168.960 307.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 336.040 1168.960 337.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 366.040 1168.960 367.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.040 1168.960 397.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 426.040 1168.960 427.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 456.040 1168.960 457.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 486.040 1168.960 487.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 516.040 1168.960 517.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.040 1168.960 547.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 576.040 1168.960 577.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 606.040 1168.960 607.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.040 1168.960 637.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 666.040 1168.960 667.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.040 1168.960 697.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 726.040 1168.960 727.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 756.040 1168.960 757.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.040 1168.960 787.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.040 1168.960 817.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.040 1168.960 847.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 876.040 1168.960 877.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 906.040 1168.960 907.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 936.040 1168.960 937.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 966.040 1168.960 967.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.040 1168.960 997.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1026.040 1168.960 1027.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.040 10.640 37.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.040 10.640 67.640 1588.720 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 81.040 371.460 82.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.040 371.460 112.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 371.460 142.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 371.460 172.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 371.460 202.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 371.460 232.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 371.460 262.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 371.460 292.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 371.460 322.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 371.460 352.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 371.460 382.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 371.460 412.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 371.460 442.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 371.460 472.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 371.460 502.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 371.460 532.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.040 371.460 562.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.040 371.460 592.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 371.460 622.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 651.040 371.460 652.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 681.040 371.460 682.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.040 371.460 712.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 371.460 742.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 371.460 772.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.040 371.460 802.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.040 371.460 832.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 861.040 371.460 862.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 891.040 371.460 892.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 371.460 922.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.040 371.460 952.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 981.040 371.460 982.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.040 371.460 1012.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1041.040 371.460 1042.640 431.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 1168.960 82.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.040 1168.960 112.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 1168.960 142.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 1168.960 172.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 1168.960 202.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 1168.960 232.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 1168.960 262.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 1168.960 292.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 1168.960 322.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 1168.960 352.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 1168.960 382.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 1168.960 412.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 1168.960 442.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 1168.960 472.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 1168.960 502.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 1168.960 532.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.040 1168.960 562.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.040 1168.960 592.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 1168.960 622.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 651.040 1168.960 652.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 681.040 1168.960 682.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.040 1168.960 712.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 1168.960 742.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 1168.960 772.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.040 1168.960 802.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.040 1168.960 832.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 861.040 1168.960 862.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 891.040 1168.960 892.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 1168.960 922.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.040 1168.960 952.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 981.040 1168.960 982.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.040 1168.960 1012.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1041.040 1168.960 1042.640 1228.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 1588.720 ;
    END
  END VPWR
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END addr[0]
  PIN addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END addr[10]
  PIN addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END addr[11]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END addr[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END clk
  PIN clk_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END clk_en
  PIN read_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END read_data[0]
  PIN read_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 742.600 4.000 743.200 ;
    END
  END read_data[10]
  PIN read_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 753.480 4.000 754.080 ;
    END
  END read_data[11]
  PIN read_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END read_data[12]
  PIN read_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END read_data[13]
  PIN read_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 787.480 4.000 788.080 ;
    END
  END read_data[14]
  PIN read_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END read_data[15]
  PIN read_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 810.600 4.000 811.200 ;
    END
  END read_data[16]
  PIN read_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.160 4.000 822.760 ;
    END
  END read_data[17]
  PIN read_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END read_data[18]
  PIN read_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 844.600 4.000 845.200 ;
    END
  END read_data[19]
  PIN read_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END read_data[1]
  PIN read_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.160 4.000 856.760 ;
    END
  END read_data[20]
  PIN read_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END read_data[21]
  PIN read_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 878.600 4.000 879.200 ;
    END
  END read_data[22]
  PIN read_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.160 4.000 890.760 ;
    END
  END read_data[23]
  PIN read_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.040 4.000 901.640 ;
    END
  END read_data[24]
  PIN read_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 912.600 4.000 913.200 ;
    END
  END read_data[25]
  PIN read_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.160 4.000 924.760 ;
    END
  END read_data[26]
  PIN read_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 935.040 4.000 935.640 ;
    END
  END read_data[27]
  PIN read_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 946.600 4.000 947.200 ;
    END
  END read_data[28]
  PIN read_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.160 4.000 958.760 ;
    END
  END read_data[29]
  PIN read_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 651.480 4.000 652.080 ;
    END
  END read_data[2]
  PIN read_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END read_data[30]
  PIN read_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END read_data[31]
  PIN read_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.160 4.000 992.760 ;
    END
  END read_data[32]
  PIN read_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END read_data[33]
  PIN read_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1014.600 4.000 1015.200 ;
    END
  END read_data[34]
  PIN read_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.160 4.000 1026.760 ;
    END
  END read_data[35]
  PIN read_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.040 4.000 1037.640 ;
    END
  END read_data[36]
  PIN read_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1048.600 4.000 1049.200 ;
    END
  END read_data[37]
  PIN read_data[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.160 4.000 1060.760 ;
    END
  END read_data[38]
  PIN read_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END read_data[3]
  PIN read_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END read_data[4]
  PIN read_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END read_data[5]
  PIN read_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END read_data[6]
  PIN read_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END read_data[7]
  PIN read_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END read_data[8]
  PIN read_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END read_data[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END rst
  PIN write_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END write_data[0]
  PIN write_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END write_data[10]
  PIN write_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END write_data[11]
  PIN write_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END write_data[12]
  PIN write_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END write_data[13]
  PIN write_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END write_data[14]
  PIN write_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END write_data[15]
  PIN write_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END write_data[16]
  PIN write_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END write_data[17]
  PIN write_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END write_data[18]
  PIN write_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END write_data[19]
  PIN write_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END write_data[1]
  PIN write_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END write_data[20]
  PIN write_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END write_data[21]
  PIN write_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.920 4.000 436.520 ;
    END
  END write_data[22]
  PIN write_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END write_data[23]
  PIN write_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END write_data[24]
  PIN write_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.920 4.000 470.520 ;
    END
  END write_data[25]
  PIN write_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END write_data[26]
  PIN write_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END write_data[27]
  PIN write_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.920 4.000 504.520 ;
    END
  END write_data[28]
  PIN write_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END write_data[29]
  PIN write_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END write_data[2]
  PIN write_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END write_data[30]
  PIN write_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END write_data[31]
  PIN write_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END write_data[32]
  PIN write_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END write_data[33]
  PIN write_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END write_data[34]
  PIN write_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END write_data[35]
  PIN write_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END write_data[36]
  PIN write_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END write_data[37]
  PIN write_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END write_data[38]
  PIN write_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END write_data[3]
  PIN write_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END write_data[4]
  PIN write_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END write_data[5]
  PIN write_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END write_data[6]
  PIN write_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END write_data[7]
  PIN write_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END write_data[8]
  PIN write_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END write_data[9]
  PIN write_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END write_en
  OBS
      LAYER li1 ;
        RECT 5.520 1167.475 1050.000 1588.565 ;
        RECT 5.520 450.245 1050.035 1167.475 ;
        RECT 5.520 447.695 1050.000 450.245 ;
        RECT 5.520 414.545 1050.035 447.695 ;
        RECT 5.520 10.795 1050.000 414.545 ;
      LAYER met1 ;
        RECT 5.520 449.380 1050.000 1594.380 ;
        RECT 5.520 446.520 1050.020 449.380 ;
        RECT 5.520 5.620 1050.000 446.520 ;
      LAYER met2 ;
        RECT 6.990 1193.770 1050.000 1594.380 ;
        RECT 6.990 275.930 1050.020 1193.770 ;
        RECT 6.990 5.595 1050.000 275.930 ;
      LAYER met3 ;
        RECT 4.000 1061.160 1049.655 1595.000 ;
        RECT 4.400 1059.760 1049.655 1061.160 ;
        RECT 4.000 1049.600 1049.655 1059.760 ;
        RECT 4.400 1048.200 1049.655 1049.600 ;
        RECT 4.000 1038.040 1049.655 1048.200 ;
        RECT 4.400 1036.640 1049.655 1038.040 ;
        RECT 4.000 1027.160 1049.655 1036.640 ;
        RECT 4.400 1025.760 1049.655 1027.160 ;
        RECT 4.000 1015.600 1049.655 1025.760 ;
        RECT 4.400 1014.200 1049.655 1015.600 ;
        RECT 4.000 1004.040 1049.655 1014.200 ;
        RECT 4.400 1002.640 1049.655 1004.040 ;
        RECT 4.000 993.160 1049.655 1002.640 ;
        RECT 4.400 991.760 1049.655 993.160 ;
        RECT 4.000 981.600 1049.655 991.760 ;
        RECT 4.400 980.200 1049.655 981.600 ;
        RECT 4.000 970.040 1049.655 980.200 ;
        RECT 4.400 968.640 1049.655 970.040 ;
        RECT 4.000 959.160 1049.655 968.640 ;
        RECT 4.400 957.760 1049.655 959.160 ;
        RECT 4.000 947.600 1049.655 957.760 ;
        RECT 4.400 946.200 1049.655 947.600 ;
        RECT 4.000 936.040 1049.655 946.200 ;
        RECT 4.400 934.640 1049.655 936.040 ;
        RECT 4.000 925.160 1049.655 934.640 ;
        RECT 4.400 923.760 1049.655 925.160 ;
        RECT 4.000 913.600 1049.655 923.760 ;
        RECT 4.400 912.200 1049.655 913.600 ;
        RECT 4.000 902.040 1049.655 912.200 ;
        RECT 4.400 900.640 1049.655 902.040 ;
        RECT 4.000 891.160 1049.655 900.640 ;
        RECT 4.400 889.760 1049.655 891.160 ;
        RECT 4.000 879.600 1049.655 889.760 ;
        RECT 4.400 878.200 1049.655 879.600 ;
        RECT 4.000 868.040 1049.655 878.200 ;
        RECT 4.400 866.640 1049.655 868.040 ;
        RECT 4.000 857.160 1049.655 866.640 ;
        RECT 4.400 855.760 1049.655 857.160 ;
        RECT 4.000 845.600 1049.655 855.760 ;
        RECT 4.400 844.200 1049.655 845.600 ;
        RECT 4.000 834.040 1049.655 844.200 ;
        RECT 4.400 832.640 1049.655 834.040 ;
        RECT 4.000 823.160 1049.655 832.640 ;
        RECT 4.400 821.760 1049.655 823.160 ;
        RECT 4.000 811.600 1049.655 821.760 ;
        RECT 4.400 810.200 1049.655 811.600 ;
        RECT 4.000 800.040 1049.655 810.200 ;
        RECT 4.400 798.640 1049.655 800.040 ;
        RECT 4.000 788.480 1049.655 798.640 ;
        RECT 4.400 787.080 1049.655 788.480 ;
        RECT 4.000 777.600 1049.655 787.080 ;
        RECT 4.400 776.200 1049.655 777.600 ;
        RECT 4.000 766.040 1049.655 776.200 ;
        RECT 4.400 764.640 1049.655 766.040 ;
        RECT 4.000 754.480 1049.655 764.640 ;
        RECT 4.400 753.080 1049.655 754.480 ;
        RECT 4.000 743.600 1049.655 753.080 ;
        RECT 4.400 742.200 1049.655 743.600 ;
        RECT 4.000 732.040 1049.655 742.200 ;
        RECT 4.400 730.640 1049.655 732.040 ;
        RECT 4.000 720.480 1049.655 730.640 ;
        RECT 4.400 719.080 1049.655 720.480 ;
        RECT 4.000 709.600 1049.655 719.080 ;
        RECT 4.400 708.200 1049.655 709.600 ;
        RECT 4.000 698.040 1049.655 708.200 ;
        RECT 4.400 696.640 1049.655 698.040 ;
        RECT 4.000 686.480 1049.655 696.640 ;
        RECT 4.400 685.080 1049.655 686.480 ;
        RECT 4.000 675.600 1049.655 685.080 ;
        RECT 4.400 674.200 1049.655 675.600 ;
        RECT 4.000 664.040 1049.655 674.200 ;
        RECT 4.400 662.640 1049.655 664.040 ;
        RECT 4.000 652.480 1049.655 662.640 ;
        RECT 4.400 651.080 1049.655 652.480 ;
        RECT 4.000 641.600 1049.655 651.080 ;
        RECT 4.400 640.200 1049.655 641.600 ;
        RECT 4.000 630.040 1049.655 640.200 ;
        RECT 4.400 628.640 1049.655 630.040 ;
        RECT 4.000 618.480 1049.655 628.640 ;
        RECT 4.400 617.080 1049.655 618.480 ;
        RECT 4.000 607.600 1049.655 617.080 ;
        RECT 4.400 606.200 1049.655 607.600 ;
        RECT 4.000 596.040 1049.655 606.200 ;
        RECT 4.400 594.640 1049.655 596.040 ;
        RECT 4.000 584.480 1049.655 594.640 ;
        RECT 4.400 583.080 1049.655 584.480 ;
        RECT 4.000 573.600 1049.655 583.080 ;
        RECT 4.400 572.200 1049.655 573.600 ;
        RECT 4.000 562.040 1049.655 572.200 ;
        RECT 4.400 560.640 1049.655 562.040 ;
        RECT 4.000 550.480 1049.655 560.640 ;
        RECT 4.400 549.080 1049.655 550.480 ;
        RECT 4.000 539.600 1049.655 549.080 ;
        RECT 4.400 538.200 1049.655 539.600 ;
        RECT 4.000 528.040 1049.655 538.200 ;
        RECT 4.400 526.640 1049.655 528.040 ;
        RECT 4.000 516.480 1049.655 526.640 ;
        RECT 4.400 515.080 1049.655 516.480 ;
        RECT 4.000 504.920 1049.655 515.080 ;
        RECT 4.400 503.520 1049.655 504.920 ;
        RECT 4.000 494.040 1049.655 503.520 ;
        RECT 4.400 492.640 1049.655 494.040 ;
        RECT 4.000 482.480 1049.655 492.640 ;
        RECT 4.400 481.080 1049.655 482.480 ;
        RECT 4.000 470.920 1049.655 481.080 ;
        RECT 4.400 469.520 1049.655 470.920 ;
        RECT 4.000 460.040 1049.655 469.520 ;
        RECT 4.400 458.640 1049.655 460.040 ;
        RECT 4.000 448.480 1049.655 458.640 ;
        RECT 4.400 447.080 1049.655 448.480 ;
        RECT 4.000 436.920 1049.655 447.080 ;
        RECT 4.400 435.520 1049.655 436.920 ;
        RECT 4.000 426.040 1049.655 435.520 ;
        RECT 4.400 424.640 1049.655 426.040 ;
        RECT 4.000 414.480 1049.655 424.640 ;
        RECT 4.400 413.080 1049.655 414.480 ;
        RECT 4.000 402.920 1049.655 413.080 ;
        RECT 4.400 401.520 1049.655 402.920 ;
        RECT 4.000 392.040 1049.655 401.520 ;
        RECT 4.400 390.640 1049.655 392.040 ;
        RECT 4.000 380.480 1049.655 390.640 ;
        RECT 4.400 379.080 1049.655 380.480 ;
        RECT 4.000 368.920 1049.655 379.080 ;
        RECT 4.400 367.520 1049.655 368.920 ;
        RECT 4.000 358.040 1049.655 367.520 ;
        RECT 4.400 356.640 1049.655 358.040 ;
        RECT 4.000 346.480 1049.655 356.640 ;
        RECT 4.400 345.080 1049.655 346.480 ;
        RECT 4.000 334.920 1049.655 345.080 ;
        RECT 4.400 333.520 1049.655 334.920 ;
        RECT 4.000 324.040 1049.655 333.520 ;
        RECT 4.400 322.640 1049.655 324.040 ;
        RECT 4.000 312.480 1049.655 322.640 ;
        RECT 4.400 311.080 1049.655 312.480 ;
        RECT 4.000 300.920 1049.655 311.080 ;
        RECT 4.400 299.520 1049.655 300.920 ;
        RECT 4.000 290.040 1049.655 299.520 ;
        RECT 4.400 288.640 1049.655 290.040 ;
        RECT 4.000 278.480 1049.655 288.640 ;
        RECT 4.400 277.080 1049.655 278.480 ;
        RECT 4.000 266.920 1049.655 277.080 ;
        RECT 4.400 265.520 1049.655 266.920 ;
        RECT 4.000 255.360 1049.655 265.520 ;
        RECT 4.400 253.960 1049.655 255.360 ;
        RECT 4.000 244.480 1049.655 253.960 ;
        RECT 4.400 243.080 1049.655 244.480 ;
        RECT 4.000 232.920 1049.655 243.080 ;
        RECT 4.400 231.520 1049.655 232.920 ;
        RECT 4.000 221.360 1049.655 231.520 ;
        RECT 4.400 219.960 1049.655 221.360 ;
        RECT 4.000 210.480 1049.655 219.960 ;
        RECT 4.400 209.080 1049.655 210.480 ;
        RECT 4.000 198.920 1049.655 209.080 ;
        RECT 4.400 197.520 1049.655 198.920 ;
        RECT 4.000 187.360 1049.655 197.520 ;
        RECT 4.400 185.960 1049.655 187.360 ;
        RECT 4.000 176.480 1049.655 185.960 ;
        RECT 4.400 175.080 1049.655 176.480 ;
        RECT 4.000 164.920 1049.655 175.080 ;
        RECT 4.400 163.520 1049.655 164.920 ;
        RECT 4.000 153.360 1049.655 163.520 ;
        RECT 4.400 151.960 1049.655 153.360 ;
        RECT 4.000 142.480 1049.655 151.960 ;
        RECT 4.400 141.080 1049.655 142.480 ;
        RECT 4.000 130.920 1049.655 141.080 ;
        RECT 4.400 129.520 1049.655 130.920 ;
        RECT 4.000 119.360 1049.655 129.520 ;
        RECT 4.400 117.960 1049.655 119.360 ;
        RECT 4.000 108.480 1049.655 117.960 ;
        RECT 4.400 107.080 1049.655 108.480 ;
        RECT 4.000 96.920 1049.655 107.080 ;
        RECT 4.400 95.520 1049.655 96.920 ;
        RECT 4.000 85.360 1049.655 95.520 ;
        RECT 4.400 83.960 1049.655 85.360 ;
        RECT 4.000 74.480 1049.655 83.960 ;
        RECT 4.400 73.080 1049.655 74.480 ;
        RECT 4.000 62.920 1049.655 73.080 ;
        RECT 4.400 61.520 1049.655 62.920 ;
        RECT 4.000 51.360 1049.655 61.520 ;
        RECT 4.400 49.960 1049.655 51.360 ;
        RECT 4.000 40.480 1049.655 49.960 ;
        RECT 4.400 39.080 1049.655 40.480 ;
        RECT 4.000 28.920 1049.655 39.080 ;
        RECT 4.400 27.520 1049.655 28.920 ;
        RECT 4.000 17.360 1049.655 27.520 ;
        RECT 4.400 15.960 1049.655 17.360 ;
        RECT 4.000 6.480 1049.655 15.960 ;
        RECT 4.400 5.080 1049.655 6.480 ;
        RECT 4.000 5.000 1049.655 5.080 ;
      LAYER met4 ;
        RECT 8.150 1589.120 1046.665 1595.000 ;
        RECT 8.150 10.240 20.640 1589.120 ;
        RECT 23.040 10.240 35.640 1589.120 ;
        RECT 38.040 10.240 50.640 1589.120 ;
        RECT 53.040 10.240 65.640 1589.120 ;
        RECT 68.040 1228.940 1046.665 1589.120 ;
        RECT 68.040 1168.560 80.640 1228.940 ;
        RECT 83.040 1168.560 95.640 1228.940 ;
        RECT 98.040 1168.560 110.640 1228.940 ;
        RECT 113.040 1168.560 125.640 1228.940 ;
        RECT 128.040 1168.560 140.640 1228.940 ;
        RECT 143.040 1168.560 155.640 1228.940 ;
        RECT 158.040 1168.560 170.640 1228.940 ;
        RECT 173.040 1168.560 185.640 1228.940 ;
        RECT 188.040 1168.560 200.640 1228.940 ;
        RECT 203.040 1168.560 215.640 1228.940 ;
        RECT 218.040 1168.560 230.640 1228.940 ;
        RECT 233.040 1168.560 245.640 1228.940 ;
        RECT 248.040 1168.560 260.640 1228.940 ;
        RECT 263.040 1168.560 275.640 1228.940 ;
        RECT 278.040 1168.560 290.640 1228.940 ;
        RECT 293.040 1168.560 305.640 1228.940 ;
        RECT 308.040 1168.560 320.640 1228.940 ;
        RECT 323.040 1168.560 335.640 1228.940 ;
        RECT 338.040 1168.560 350.640 1228.940 ;
        RECT 353.040 1168.560 365.640 1228.940 ;
        RECT 368.040 1168.560 380.640 1228.940 ;
        RECT 383.040 1168.560 395.640 1228.940 ;
        RECT 398.040 1168.560 410.640 1228.940 ;
        RECT 413.040 1168.560 425.640 1228.940 ;
        RECT 428.040 1168.560 440.640 1228.940 ;
        RECT 443.040 1168.560 455.640 1228.940 ;
        RECT 458.040 1168.560 470.640 1228.940 ;
        RECT 473.040 1168.560 485.640 1228.940 ;
        RECT 488.040 1168.560 500.640 1228.940 ;
        RECT 503.040 1168.560 515.640 1228.940 ;
        RECT 518.040 1168.560 530.640 1228.940 ;
        RECT 533.040 1168.560 545.640 1228.940 ;
        RECT 548.040 1168.560 560.640 1228.940 ;
        RECT 563.040 1168.560 575.640 1228.940 ;
        RECT 578.040 1168.560 590.640 1228.940 ;
        RECT 593.040 1168.560 605.640 1228.940 ;
        RECT 608.040 1168.560 620.640 1228.940 ;
        RECT 623.040 1168.560 635.640 1228.940 ;
        RECT 638.040 1168.560 650.640 1228.940 ;
        RECT 653.040 1168.560 665.640 1228.940 ;
        RECT 668.040 1168.560 680.640 1228.940 ;
        RECT 683.040 1168.560 695.640 1228.940 ;
        RECT 698.040 1168.560 710.640 1228.940 ;
        RECT 713.040 1168.560 725.640 1228.940 ;
        RECT 728.040 1168.560 740.640 1228.940 ;
        RECT 743.040 1168.560 755.640 1228.940 ;
        RECT 758.040 1168.560 770.640 1228.940 ;
        RECT 773.040 1168.560 785.640 1228.940 ;
        RECT 788.040 1168.560 800.640 1228.940 ;
        RECT 803.040 1168.560 815.640 1228.940 ;
        RECT 818.040 1168.560 830.640 1228.940 ;
        RECT 833.040 1168.560 845.640 1228.940 ;
        RECT 848.040 1168.560 860.640 1228.940 ;
        RECT 863.040 1168.560 875.640 1228.940 ;
        RECT 878.040 1168.560 890.640 1228.940 ;
        RECT 893.040 1168.560 905.640 1228.940 ;
        RECT 908.040 1168.560 920.640 1228.940 ;
        RECT 923.040 1168.560 935.640 1228.940 ;
        RECT 938.040 1168.560 950.640 1228.940 ;
        RECT 953.040 1168.560 965.640 1228.940 ;
        RECT 968.040 1168.560 980.640 1228.940 ;
        RECT 983.040 1168.560 995.640 1228.940 ;
        RECT 998.040 1168.560 1010.640 1228.940 ;
        RECT 1013.040 1168.560 1025.640 1228.940 ;
        RECT 1028.040 1168.560 1040.640 1228.940 ;
        RECT 1043.040 1168.560 1046.665 1228.940 ;
        RECT 68.040 431.440 1046.665 1168.560 ;
        RECT 68.040 371.060 80.640 431.440 ;
        RECT 83.040 371.060 95.640 431.440 ;
        RECT 98.040 371.060 110.640 431.440 ;
        RECT 113.040 371.060 125.640 431.440 ;
        RECT 128.040 371.060 140.640 431.440 ;
        RECT 143.040 371.060 155.640 431.440 ;
        RECT 158.040 371.060 170.640 431.440 ;
        RECT 173.040 371.060 185.640 431.440 ;
        RECT 188.040 371.060 200.640 431.440 ;
        RECT 203.040 371.060 215.640 431.440 ;
        RECT 218.040 371.060 230.640 431.440 ;
        RECT 233.040 371.060 245.640 431.440 ;
        RECT 248.040 371.060 260.640 431.440 ;
        RECT 263.040 371.060 275.640 431.440 ;
        RECT 278.040 371.060 290.640 431.440 ;
        RECT 293.040 371.060 305.640 431.440 ;
        RECT 308.040 371.060 320.640 431.440 ;
        RECT 323.040 371.060 335.640 431.440 ;
        RECT 338.040 371.060 350.640 431.440 ;
        RECT 353.040 371.060 365.640 431.440 ;
        RECT 368.040 371.060 380.640 431.440 ;
        RECT 383.040 371.060 395.640 431.440 ;
        RECT 398.040 371.060 410.640 431.440 ;
        RECT 413.040 371.060 425.640 431.440 ;
        RECT 428.040 371.060 440.640 431.440 ;
        RECT 443.040 371.060 455.640 431.440 ;
        RECT 458.040 371.060 470.640 431.440 ;
        RECT 473.040 371.060 485.640 431.440 ;
        RECT 488.040 371.060 500.640 431.440 ;
        RECT 503.040 371.060 515.640 431.440 ;
        RECT 518.040 371.060 530.640 431.440 ;
        RECT 533.040 371.060 545.640 431.440 ;
        RECT 548.040 371.060 560.640 431.440 ;
        RECT 563.040 371.060 575.640 431.440 ;
        RECT 578.040 371.060 590.640 431.440 ;
        RECT 593.040 371.060 605.640 431.440 ;
        RECT 608.040 371.060 620.640 431.440 ;
        RECT 623.040 371.060 635.640 431.440 ;
        RECT 638.040 371.060 650.640 431.440 ;
        RECT 653.040 371.060 665.640 431.440 ;
        RECT 668.040 371.060 680.640 431.440 ;
        RECT 683.040 371.060 695.640 431.440 ;
        RECT 698.040 371.060 710.640 431.440 ;
        RECT 713.040 371.060 725.640 431.440 ;
        RECT 728.040 371.060 740.640 431.440 ;
        RECT 743.040 371.060 755.640 431.440 ;
        RECT 758.040 371.060 770.640 431.440 ;
        RECT 773.040 371.060 785.640 431.440 ;
        RECT 788.040 371.060 800.640 431.440 ;
        RECT 803.040 371.060 815.640 431.440 ;
        RECT 818.040 371.060 830.640 431.440 ;
        RECT 833.040 371.060 845.640 431.440 ;
        RECT 848.040 371.060 860.640 431.440 ;
        RECT 863.040 371.060 875.640 431.440 ;
        RECT 878.040 371.060 890.640 431.440 ;
        RECT 893.040 371.060 905.640 431.440 ;
        RECT 908.040 371.060 920.640 431.440 ;
        RECT 923.040 371.060 935.640 431.440 ;
        RECT 938.040 371.060 950.640 431.440 ;
        RECT 953.040 371.060 965.640 431.440 ;
        RECT 968.040 371.060 980.640 431.440 ;
        RECT 983.040 371.060 995.640 431.440 ;
        RECT 998.040 371.060 1010.640 431.440 ;
        RECT 1013.040 371.060 1025.640 431.440 ;
        RECT 1028.040 371.060 1040.640 431.440 ;
        RECT 1043.040 371.060 1046.665 431.440 ;
        RECT 68.040 10.240 1046.665 371.060 ;
        RECT 8.150 5.000 1046.665 10.240 ;
      LAYER met5 ;
        RECT 7.940 436.100 815.460 1178.900 ;
  END
END sram_39_4096
END LIBRARY

