VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sram_32_4096
  CLASS BLOCK ;
  FOREIGN sram_32_4096 ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 1600.000 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.040 365.340 97.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.040 365.340 127.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 156.040 365.340 157.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 186.040 365.340 187.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 216.040 365.340 217.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.040 365.340 247.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 276.040 365.340 277.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 306.040 365.340 307.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 336.040 365.340 337.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 366.040 365.340 367.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.040 365.340 397.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 426.040 365.340 427.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 456.040 365.340 457.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 486.040 365.340 487.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 516.040 365.340 517.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.040 365.340 547.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 576.040 365.340 577.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 606.040 365.340 607.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.040 365.340 637.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 666.040 365.340 667.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.040 365.340 697.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 726.040 365.340 727.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 756.040 365.340 757.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.040 365.340 787.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.040 365.340 817.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.040 365.340 847.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 876.040 365.340 877.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.040 1162.840 97.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.040 1162.840 127.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 156.040 1162.840 157.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 186.040 1162.840 187.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 216.040 1162.840 217.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.040 1162.840 247.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 276.040 1162.840 277.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 306.040 1162.840 307.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 336.040 1162.840 337.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 366.040 1162.840 367.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.040 1162.840 397.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 426.040 1162.840 427.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 456.040 1162.840 457.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 486.040 1162.840 487.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 516.040 1162.840 517.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.040 1162.840 547.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 576.040 1162.840 577.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 606.040 1162.840 607.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.040 1162.840 637.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 666.040 1162.840 667.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.040 1162.840 697.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 726.040 1162.840 727.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 756.040 1162.840 757.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.040 1162.840 787.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.040 1162.840 817.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.040 1162.840 847.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 876.040 1162.840 877.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.040 10.640 37.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.040 10.640 67.640 1588.720 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 81.040 365.340 82.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.040 365.340 112.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 365.340 142.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 365.340 172.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 365.340 202.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 365.340 232.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 365.340 262.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 365.340 292.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 365.340 322.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 365.340 352.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 365.340 382.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 365.340 412.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 365.340 442.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 365.340 472.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 365.340 502.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 365.340 532.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.040 365.340 562.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.040 365.340 592.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 365.340 622.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 651.040 365.340 652.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 681.040 365.340 682.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.040 365.340 712.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 365.340 742.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 365.340 772.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.040 365.340 802.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.040 365.340 832.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 861.040 365.340 862.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 891.040 365.340 892.640 437.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 1162.840 82.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.040 1162.840 112.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 1162.840 142.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 1162.840 172.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 1162.840 202.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 1162.840 232.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 1162.840 262.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 1162.840 292.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 1162.840 322.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 1162.840 352.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 1162.840 382.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 1162.840 412.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 1162.840 442.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 1162.840 472.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 1162.840 502.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 1162.840 532.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.040 1162.840 562.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.040 1162.840 592.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 1162.840 622.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 651.040 1162.840 652.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 681.040 1162.840 682.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.040 1162.840 712.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 1162.840 742.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 1162.840 772.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.040 1162.840 802.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.040 1162.840 832.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 861.040 1162.840 862.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 891.040 1162.840 892.640 1234.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 1588.720 ;
    END
  END VPWR
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END addr[0]
  PIN addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END addr[10]
  PIN addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END addr[11]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END addr[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END clk
  PIN clk_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END clk_en
  PIN read_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 645.360 4.000 645.960 ;
    END
  END read_data[0]
  PIN read_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END read_data[10]
  PIN read_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END read_data[11]
  PIN read_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END read_data[12]
  PIN read_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.760 4.000 819.360 ;
    END
  END read_data[13]
  PIN read_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END read_data[14]
  PIN read_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.280 4.000 845.880 ;
    END
  END read_data[15]
  PIN read_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.880 4.000 859.480 ;
    END
  END read_data[16]
  PIN read_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 872.480 4.000 873.080 ;
    END
  END read_data[17]
  PIN read_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 885.400 4.000 886.000 ;
    END
  END read_data[18]
  PIN read_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.000 4.000 899.600 ;
    END
  END read_data[19]
  PIN read_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.960 4.000 659.560 ;
    END
  END read_data[1]
  PIN read_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.920 4.000 912.520 ;
    END
  END read_data[20]
  PIN read_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 925.520 4.000 926.120 ;
    END
  END read_data[21]
  PIN read_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.120 4.000 939.720 ;
    END
  END read_data[22]
  PIN read_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END read_data[23]
  PIN read_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END read_data[24]
  PIN read_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 978.560 4.000 979.160 ;
    END
  END read_data[25]
  PIN read_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.160 4.000 992.760 ;
    END
  END read_data[26]
  PIN read_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1005.760 4.000 1006.360 ;
    END
  END read_data[27]
  PIN read_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.680 4.000 1019.280 ;
    END
  END read_data[28]
  PIN read_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.280 4.000 1032.880 ;
    END
  END read_data[29]
  PIN read_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 672.560 4.000 673.160 ;
    END
  END read_data[2]
  PIN read_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1045.200 4.000 1045.800 ;
    END
  END read_data[30]
  PIN read_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1058.800 4.000 1059.400 ;
    END
  END read_data[31]
  PIN read_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END read_data[3]
  PIN read_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END read_data[4]
  PIN read_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.000 4.000 712.600 ;
    END
  END read_data[5]
  PIN read_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 725.600 4.000 726.200 ;
    END
  END read_data[6]
  PIN read_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.200 4.000 739.800 ;
    END
  END read_data[7]
  PIN read_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END read_data[8]
  PIN read_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.720 4.000 766.320 ;
    END
  END read_data[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END rst
  PIN write_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END write_data[0]
  PIN write_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END write_data[10]
  PIN write_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END write_data[11]
  PIN write_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END write_data[12]
  PIN write_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END write_data[13]
  PIN write_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.000 4.000 406.600 ;
    END
  END write_data[14]
  PIN write_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END write_data[15]
  PIN write_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END write_data[16]
  PIN write_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END write_data[17]
  PIN write_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END write_data[18]
  PIN write_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END write_data[19]
  PIN write_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END write_data[1]
  PIN write_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END write_data[20]
  PIN write_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END write_data[21]
  PIN write_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.080 4.000 512.680 ;
    END
  END write_data[22]
  PIN write_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.680 4.000 526.280 ;
    END
  END write_data[23]
  PIN write_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.280 4.000 539.880 ;
    END
  END write_data[24]
  PIN write_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END write_data[25]
  PIN write_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END write_data[26]
  PIN write_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END write_data[27]
  PIN write_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 592.320 4.000 592.920 ;
    END
  END write_data[28]
  PIN write_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.920 4.000 606.520 ;
    END
  END write_data[29]
  PIN write_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END write_data[2]
  PIN write_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END write_data[30]
  PIN write_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END write_data[31]
  PIN write_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END write_data[3]
  PIN write_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.720 4.000 273.320 ;
    END
  END write_data[4]
  PIN write_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END write_data[5]
  PIN write_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END write_data[6]
  PIN write_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END write_data[7]
  PIN write_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END write_data[8]
  PIN write_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END write_data[9]
  PIN write_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END write_en
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 1588.565 ;
      LAYER met1 ;
        RECT 5.520 1128.020 900.000 1594.380 ;
        RECT 5.520 1124.140 900.060 1128.020 ;
        RECT 5.520 449.720 900.000 1124.140 ;
        RECT 5.520 447.880 900.060 449.720 ;
        RECT 5.520 5.620 900.000 447.880 ;
      LAYER met2 ;
        RECT 6.990 1167.290 900.000 1594.380 ;
        RECT 6.990 1126.350 900.060 1167.290 ;
        RECT 6.990 1125.300 900.000 1126.350 ;
        RECT 6.990 449.750 900.060 1125.300 ;
        RECT 6.990 448.570 900.000 449.750 ;
        RECT 6.990 431.390 900.060 448.570 ;
        RECT 6.990 5.620 900.000 431.390 ;
      LAYER met3 ;
        RECT 4.000 1059.800 899.695 1595.000 ;
        RECT 4.400 1058.400 899.695 1059.800 ;
        RECT 4.000 1046.200 899.695 1058.400 ;
        RECT 4.400 1044.800 899.695 1046.200 ;
        RECT 4.000 1033.280 899.695 1044.800 ;
        RECT 4.400 1031.880 899.695 1033.280 ;
        RECT 4.000 1019.680 899.695 1031.880 ;
        RECT 4.400 1018.280 899.695 1019.680 ;
        RECT 4.000 1006.760 899.695 1018.280 ;
        RECT 4.400 1005.360 899.695 1006.760 ;
        RECT 4.000 993.160 899.695 1005.360 ;
        RECT 4.400 991.760 899.695 993.160 ;
        RECT 4.000 979.560 899.695 991.760 ;
        RECT 4.400 978.160 899.695 979.560 ;
        RECT 4.000 966.640 899.695 978.160 ;
        RECT 4.400 965.240 899.695 966.640 ;
        RECT 4.000 953.040 899.695 965.240 ;
        RECT 4.400 951.640 899.695 953.040 ;
        RECT 4.000 940.120 899.695 951.640 ;
        RECT 4.400 938.720 899.695 940.120 ;
        RECT 4.000 926.520 899.695 938.720 ;
        RECT 4.400 925.120 899.695 926.520 ;
        RECT 4.000 912.920 899.695 925.120 ;
        RECT 4.400 911.520 899.695 912.920 ;
        RECT 4.000 900.000 899.695 911.520 ;
        RECT 4.400 898.600 899.695 900.000 ;
        RECT 4.000 886.400 899.695 898.600 ;
        RECT 4.400 885.000 899.695 886.400 ;
        RECT 4.000 873.480 899.695 885.000 ;
        RECT 4.400 872.080 899.695 873.480 ;
        RECT 4.000 859.880 899.695 872.080 ;
        RECT 4.400 858.480 899.695 859.880 ;
        RECT 4.000 846.280 899.695 858.480 ;
        RECT 4.400 844.880 899.695 846.280 ;
        RECT 4.000 833.360 899.695 844.880 ;
        RECT 4.400 831.960 899.695 833.360 ;
        RECT 4.000 819.760 899.695 831.960 ;
        RECT 4.400 818.360 899.695 819.760 ;
        RECT 4.000 806.840 899.695 818.360 ;
        RECT 4.400 805.440 899.695 806.840 ;
        RECT 4.000 793.240 899.695 805.440 ;
        RECT 4.400 791.840 899.695 793.240 ;
        RECT 4.000 779.640 899.695 791.840 ;
        RECT 4.400 778.240 899.695 779.640 ;
        RECT 4.000 766.720 899.695 778.240 ;
        RECT 4.400 765.320 899.695 766.720 ;
        RECT 4.000 753.120 899.695 765.320 ;
        RECT 4.400 751.720 899.695 753.120 ;
        RECT 4.000 740.200 899.695 751.720 ;
        RECT 4.400 738.800 899.695 740.200 ;
        RECT 4.000 726.600 899.695 738.800 ;
        RECT 4.400 725.200 899.695 726.600 ;
        RECT 4.000 713.000 899.695 725.200 ;
        RECT 4.400 711.600 899.695 713.000 ;
        RECT 4.000 700.080 899.695 711.600 ;
        RECT 4.400 698.680 899.695 700.080 ;
        RECT 4.000 686.480 899.695 698.680 ;
        RECT 4.400 685.080 899.695 686.480 ;
        RECT 4.000 673.560 899.695 685.080 ;
        RECT 4.400 672.160 899.695 673.560 ;
        RECT 4.000 659.960 899.695 672.160 ;
        RECT 4.400 658.560 899.695 659.960 ;
        RECT 4.000 646.360 899.695 658.560 ;
        RECT 4.400 644.960 899.695 646.360 ;
        RECT 4.000 633.440 899.695 644.960 ;
        RECT 4.400 632.040 899.695 633.440 ;
        RECT 4.000 619.840 899.695 632.040 ;
        RECT 4.400 618.440 899.695 619.840 ;
        RECT 4.000 606.920 899.695 618.440 ;
        RECT 4.400 605.520 899.695 606.920 ;
        RECT 4.000 593.320 899.695 605.520 ;
        RECT 4.400 591.920 899.695 593.320 ;
        RECT 4.000 579.720 899.695 591.920 ;
        RECT 4.400 578.320 899.695 579.720 ;
        RECT 4.000 566.800 899.695 578.320 ;
        RECT 4.400 565.400 899.695 566.800 ;
        RECT 4.000 553.200 899.695 565.400 ;
        RECT 4.400 551.800 899.695 553.200 ;
        RECT 4.000 540.280 899.695 551.800 ;
        RECT 4.400 538.880 899.695 540.280 ;
        RECT 4.000 526.680 899.695 538.880 ;
        RECT 4.400 525.280 899.695 526.680 ;
        RECT 4.000 513.080 899.695 525.280 ;
        RECT 4.400 511.680 899.695 513.080 ;
        RECT 4.000 500.160 899.695 511.680 ;
        RECT 4.400 498.760 899.695 500.160 ;
        RECT 4.000 486.560 899.695 498.760 ;
        RECT 4.400 485.160 899.695 486.560 ;
        RECT 4.000 473.640 899.695 485.160 ;
        RECT 4.400 472.240 899.695 473.640 ;
        RECT 4.000 460.040 899.695 472.240 ;
        RECT 4.400 458.640 899.695 460.040 ;
        RECT 4.000 446.440 899.695 458.640 ;
        RECT 4.400 445.040 899.695 446.440 ;
        RECT 4.000 433.520 899.695 445.040 ;
        RECT 4.400 432.120 899.695 433.520 ;
        RECT 4.000 419.920 899.695 432.120 ;
        RECT 4.400 418.520 899.695 419.920 ;
        RECT 4.000 407.000 899.695 418.520 ;
        RECT 4.400 405.600 899.695 407.000 ;
        RECT 4.000 393.400 899.695 405.600 ;
        RECT 4.400 392.000 899.695 393.400 ;
        RECT 4.000 379.800 899.695 392.000 ;
        RECT 4.400 378.400 899.695 379.800 ;
        RECT 4.000 366.880 899.695 378.400 ;
        RECT 4.400 365.480 899.695 366.880 ;
        RECT 4.000 353.280 899.695 365.480 ;
        RECT 4.400 351.880 899.695 353.280 ;
        RECT 4.000 340.360 899.695 351.880 ;
        RECT 4.400 338.960 899.695 340.360 ;
        RECT 4.000 326.760 899.695 338.960 ;
        RECT 4.400 325.360 899.695 326.760 ;
        RECT 4.000 313.160 899.695 325.360 ;
        RECT 4.400 311.760 899.695 313.160 ;
        RECT 4.000 300.240 899.695 311.760 ;
        RECT 4.400 298.840 899.695 300.240 ;
        RECT 4.000 286.640 899.695 298.840 ;
        RECT 4.400 285.240 899.695 286.640 ;
        RECT 4.000 273.720 899.695 285.240 ;
        RECT 4.400 272.320 899.695 273.720 ;
        RECT 4.000 260.120 899.695 272.320 ;
        RECT 4.400 258.720 899.695 260.120 ;
        RECT 4.000 246.520 899.695 258.720 ;
        RECT 4.400 245.120 899.695 246.520 ;
        RECT 4.000 233.600 899.695 245.120 ;
        RECT 4.400 232.200 899.695 233.600 ;
        RECT 4.000 220.000 899.695 232.200 ;
        RECT 4.400 218.600 899.695 220.000 ;
        RECT 4.000 207.080 899.695 218.600 ;
        RECT 4.400 205.680 899.695 207.080 ;
        RECT 4.000 193.480 899.695 205.680 ;
        RECT 4.400 192.080 899.695 193.480 ;
        RECT 4.000 179.880 899.695 192.080 ;
        RECT 4.400 178.480 899.695 179.880 ;
        RECT 4.000 166.960 899.695 178.480 ;
        RECT 4.400 165.560 899.695 166.960 ;
        RECT 4.000 153.360 899.695 165.560 ;
        RECT 4.400 151.960 899.695 153.360 ;
        RECT 4.000 140.440 899.695 151.960 ;
        RECT 4.400 139.040 899.695 140.440 ;
        RECT 4.000 126.840 899.695 139.040 ;
        RECT 4.400 125.440 899.695 126.840 ;
        RECT 4.000 113.240 899.695 125.440 ;
        RECT 4.400 111.840 899.695 113.240 ;
        RECT 4.000 100.320 899.695 111.840 ;
        RECT 4.400 98.920 899.695 100.320 ;
        RECT 4.000 86.720 899.695 98.920 ;
        RECT 4.400 85.320 899.695 86.720 ;
        RECT 4.000 73.800 899.695 85.320 ;
        RECT 4.400 72.400 899.695 73.800 ;
        RECT 4.000 60.200 899.695 72.400 ;
        RECT 4.400 58.800 899.695 60.200 ;
        RECT 4.000 46.600 899.695 58.800 ;
        RECT 4.400 45.200 899.695 46.600 ;
        RECT 4.000 33.680 899.695 45.200 ;
        RECT 4.400 32.280 899.695 33.680 ;
        RECT 4.000 20.080 899.695 32.280 ;
        RECT 4.400 18.680 899.695 20.080 ;
        RECT 4.000 7.160 899.695 18.680 ;
        RECT 4.400 5.760 899.695 7.160 ;
        RECT 4.000 5.000 899.695 5.760 ;
      LAYER met4 ;
        RECT 19.615 1589.120 899.465 1595.000 ;
        RECT 19.615 10.240 20.640 1589.120 ;
        RECT 23.040 10.240 35.640 1589.120 ;
        RECT 38.040 10.240 50.640 1589.120 ;
        RECT 53.040 10.240 65.640 1589.120 ;
        RECT 68.040 1235.060 899.465 1589.120 ;
        RECT 68.040 1162.440 80.640 1235.060 ;
        RECT 83.040 1162.440 95.640 1235.060 ;
        RECT 98.040 1162.440 110.640 1235.060 ;
        RECT 113.040 1162.440 125.640 1235.060 ;
        RECT 128.040 1162.440 140.640 1235.060 ;
        RECT 143.040 1162.440 155.640 1235.060 ;
        RECT 158.040 1162.440 170.640 1235.060 ;
        RECT 173.040 1162.440 185.640 1235.060 ;
        RECT 188.040 1162.440 200.640 1235.060 ;
        RECT 203.040 1162.440 215.640 1235.060 ;
        RECT 218.040 1162.440 230.640 1235.060 ;
        RECT 233.040 1162.440 245.640 1235.060 ;
        RECT 248.040 1162.440 260.640 1235.060 ;
        RECT 263.040 1162.440 275.640 1235.060 ;
        RECT 278.040 1162.440 290.640 1235.060 ;
        RECT 293.040 1162.440 305.640 1235.060 ;
        RECT 308.040 1162.440 320.640 1235.060 ;
        RECT 323.040 1162.440 335.640 1235.060 ;
        RECT 338.040 1162.440 350.640 1235.060 ;
        RECT 353.040 1162.440 365.640 1235.060 ;
        RECT 368.040 1162.440 380.640 1235.060 ;
        RECT 383.040 1162.440 395.640 1235.060 ;
        RECT 398.040 1162.440 410.640 1235.060 ;
        RECT 413.040 1162.440 425.640 1235.060 ;
        RECT 428.040 1162.440 440.640 1235.060 ;
        RECT 443.040 1162.440 455.640 1235.060 ;
        RECT 458.040 1162.440 470.640 1235.060 ;
        RECT 473.040 1162.440 485.640 1235.060 ;
        RECT 488.040 1162.440 500.640 1235.060 ;
        RECT 503.040 1162.440 515.640 1235.060 ;
        RECT 518.040 1162.440 530.640 1235.060 ;
        RECT 533.040 1162.440 545.640 1235.060 ;
        RECT 548.040 1162.440 560.640 1235.060 ;
        RECT 563.040 1162.440 575.640 1235.060 ;
        RECT 578.040 1162.440 590.640 1235.060 ;
        RECT 593.040 1162.440 605.640 1235.060 ;
        RECT 608.040 1162.440 620.640 1235.060 ;
        RECT 623.040 1162.440 635.640 1235.060 ;
        RECT 638.040 1162.440 650.640 1235.060 ;
        RECT 653.040 1162.440 665.640 1235.060 ;
        RECT 668.040 1162.440 680.640 1235.060 ;
        RECT 683.040 1162.440 695.640 1235.060 ;
        RECT 698.040 1162.440 710.640 1235.060 ;
        RECT 713.040 1162.440 725.640 1235.060 ;
        RECT 728.040 1162.440 740.640 1235.060 ;
        RECT 743.040 1162.440 755.640 1235.060 ;
        RECT 758.040 1162.440 770.640 1235.060 ;
        RECT 773.040 1162.440 785.640 1235.060 ;
        RECT 788.040 1162.440 800.640 1235.060 ;
        RECT 803.040 1162.440 815.640 1235.060 ;
        RECT 818.040 1162.440 830.640 1235.060 ;
        RECT 833.040 1162.440 845.640 1235.060 ;
        RECT 848.040 1162.440 860.640 1235.060 ;
        RECT 863.040 1162.440 875.640 1235.060 ;
        RECT 878.040 1162.440 890.640 1235.060 ;
        RECT 893.040 1162.440 899.465 1235.060 ;
        RECT 68.040 437.560 899.465 1162.440 ;
        RECT 68.040 364.940 80.640 437.560 ;
        RECT 83.040 364.940 95.640 437.560 ;
        RECT 98.040 364.940 110.640 437.560 ;
        RECT 113.040 364.940 125.640 437.560 ;
        RECT 128.040 364.940 140.640 437.560 ;
        RECT 143.040 364.940 155.640 437.560 ;
        RECT 158.040 364.940 170.640 437.560 ;
        RECT 173.040 364.940 185.640 437.560 ;
        RECT 188.040 364.940 200.640 437.560 ;
        RECT 203.040 364.940 215.640 437.560 ;
        RECT 218.040 364.940 230.640 437.560 ;
        RECT 233.040 364.940 245.640 437.560 ;
        RECT 248.040 364.940 260.640 437.560 ;
        RECT 263.040 364.940 275.640 437.560 ;
        RECT 278.040 364.940 290.640 437.560 ;
        RECT 293.040 364.940 305.640 437.560 ;
        RECT 308.040 364.940 320.640 437.560 ;
        RECT 323.040 364.940 335.640 437.560 ;
        RECT 338.040 364.940 350.640 437.560 ;
        RECT 353.040 364.940 365.640 437.560 ;
        RECT 368.040 364.940 380.640 437.560 ;
        RECT 383.040 364.940 395.640 437.560 ;
        RECT 398.040 364.940 410.640 437.560 ;
        RECT 413.040 364.940 425.640 437.560 ;
        RECT 428.040 364.940 440.640 437.560 ;
        RECT 443.040 364.940 455.640 437.560 ;
        RECT 458.040 364.940 470.640 437.560 ;
        RECT 473.040 364.940 485.640 437.560 ;
        RECT 488.040 364.940 500.640 437.560 ;
        RECT 503.040 364.940 515.640 437.560 ;
        RECT 518.040 364.940 530.640 437.560 ;
        RECT 533.040 364.940 545.640 437.560 ;
        RECT 548.040 364.940 560.640 437.560 ;
        RECT 563.040 364.940 575.640 437.560 ;
        RECT 578.040 364.940 590.640 437.560 ;
        RECT 593.040 364.940 605.640 437.560 ;
        RECT 608.040 364.940 620.640 437.560 ;
        RECT 623.040 364.940 635.640 437.560 ;
        RECT 638.040 364.940 650.640 437.560 ;
        RECT 653.040 364.940 665.640 437.560 ;
        RECT 668.040 364.940 680.640 437.560 ;
        RECT 683.040 364.940 695.640 437.560 ;
        RECT 698.040 364.940 710.640 437.560 ;
        RECT 713.040 364.940 725.640 437.560 ;
        RECT 728.040 364.940 740.640 437.560 ;
        RECT 743.040 364.940 755.640 437.560 ;
        RECT 758.040 364.940 770.640 437.560 ;
        RECT 773.040 364.940 785.640 437.560 ;
        RECT 788.040 364.940 800.640 437.560 ;
        RECT 803.040 364.940 815.640 437.560 ;
        RECT 818.040 364.940 830.640 437.560 ;
        RECT 833.040 364.940 845.640 437.560 ;
        RECT 848.040 364.940 860.640 437.560 ;
        RECT 863.040 364.940 875.640 437.560 ;
        RECT 878.040 364.940 890.640 437.560 ;
        RECT 893.040 364.940 899.465 437.560 ;
        RECT 68.040 10.240 899.465 364.940 ;
        RECT 19.615 5.000 899.465 10.240 ;
      LAYER met5 ;
        RECT 76.940 1136.500 890.900 1158.500 ;
  END
END sram_32_4096
END LIBRARY

