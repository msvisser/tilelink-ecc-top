VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sram_38_4096
  CLASS BLOCK ;
  FOREIGN sram_38_4096 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1050.000 BY 1600.000 ;
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END addr[0]
  PIN addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END addr[10]
  PIN addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END addr[11]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END addr[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END clk
  PIN clk_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END clk_en
  PIN read_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END read_data[0]
  PIN read_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END read_data[10]
  PIN read_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END read_data[11]
  PIN read_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 4.000 770.400 ;
    END
  END read_data[12]
  PIN read_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 781.360 4.000 781.960 ;
    END
  END read_data[13]
  PIN read_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END read_data[14]
  PIN read_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.160 4.000 805.760 ;
    END
  END read_data[15]
  PIN read_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.720 4.000 817.320 ;
    END
  END read_data[16]
  PIN read_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END read_data[17]
  PIN read_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END read_data[18]
  PIN read_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 851.400 4.000 852.000 ;
    END
  END read_data[19]
  PIN read_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END read_data[1]
  PIN read_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.960 4.000 863.560 ;
    END
  END read_data[20]
  PIN read_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 874.520 4.000 875.120 ;
    END
  END read_data[21]
  PIN read_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.080 4.000 886.680 ;
    END
  END read_data[22]
  PIN read_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END read_data[23]
  PIN read_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.200 4.000 909.800 ;
    END
  END read_data[24]
  PIN read_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.760 4.000 921.360 ;
    END
  END read_data[25]
  PIN read_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 932.320 4.000 932.920 ;
    END
  END read_data[26]
  PIN read_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 943.880 4.000 944.480 ;
    END
  END read_data[27]
  PIN read_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END read_data[28]
  PIN read_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 967.000 4.000 967.600 ;
    END
  END read_data[29]
  PIN read_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END read_data[2]
  PIN read_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 978.560 4.000 979.160 ;
    END
  END read_data[30]
  PIN read_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.120 4.000 990.720 ;
    END
  END read_data[31]
  PIN read_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.680 4.000 1002.280 ;
    END
  END read_data[32]
  PIN read_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END read_data[33]
  PIN read_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1024.800 4.000 1025.400 ;
    END
  END read_data[34]
  PIN read_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1036.360 4.000 1036.960 ;
    END
  END read_data[35]
  PIN read_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.920 4.000 1048.520 ;
    END
  END read_data[36]
  PIN read_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1059.480 4.000 1060.080 ;
    END
  END read_data[37]
  PIN read_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.760 4.000 666.360 ;
    END
  END read_data[3]
  PIN read_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END read_data[4]
  PIN read_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.880 4.000 689.480 ;
    END
  END read_data[5]
  PIN read_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END read_data[6]
  PIN read_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.000 4.000 712.600 ;
    END
  END read_data[7]
  PIN read_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 723.560 4.000 724.160 ;
    END
  END read_data[8]
  PIN read_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.120 4.000 735.720 ;
    END
  END read_data[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 111.040 370.100 112.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 370.100 142.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 370.100 172.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 370.100 202.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 370.100 232.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 370.100 262.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 370.100 292.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 370.100 322.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 370.100 352.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 370.100 382.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 370.100 412.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 370.100 442.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 370.100 472.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 370.100 502.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 370.100 532.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.040 370.100 562.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.040 370.100 592.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 370.100 622.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 651.040 370.100 652.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 681.040 370.100 682.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.040 370.100 712.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 370.100 742.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 370.100 772.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.040 370.100 802.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.040 370.100 832.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 861.040 370.100 862.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 891.040 370.100 892.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 370.100 922.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.040 370.100 952.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 981.040 370.100 982.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.040 370.100 1012.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1041.040 370.100 1042.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.040 1167.600 112.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 1167.600 142.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 1167.600 172.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 1167.600 202.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 1167.600 232.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 1167.600 262.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 1167.600 292.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 1167.600 322.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 1167.600 352.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 1167.600 382.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 1167.600 412.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 1167.600 442.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 1167.600 472.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 1167.600 502.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 1167.600 532.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.040 1167.600 562.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.040 1167.600 592.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 1167.600 622.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 651.040 1167.600 652.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 681.040 1167.600 682.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.040 1167.600 712.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 1167.600 742.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 1167.600 772.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.040 1167.600 802.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.040 1167.600 832.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 861.040 1167.600 862.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 891.040 1167.600 892.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 1167.600 922.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.040 1167.600 952.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 981.040 1167.600 982.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.040 1167.600 1012.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1041.040 1167.600 1042.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 10.640 82.640 1588.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.040 370.100 97.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.040 370.100 127.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 156.040 370.100 157.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 186.040 370.100 187.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 216.040 370.100 217.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.040 370.100 247.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 276.040 370.100 277.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 306.040 370.100 307.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 336.040 370.100 337.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 366.040 370.100 367.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.040 370.100 397.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 426.040 370.100 427.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 456.040 370.100 457.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 486.040 370.100 487.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 516.040 370.100 517.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.040 370.100 547.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 576.040 370.100 577.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 606.040 370.100 607.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.040 370.100 637.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 666.040 370.100 667.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.040 370.100 697.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 726.040 370.100 727.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 756.040 370.100 757.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.040 370.100 787.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.040 370.100 817.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.040 370.100 847.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 876.040 370.100 877.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 906.040 370.100 907.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 936.040 370.100 937.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 966.040 370.100 967.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.040 370.100 997.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1026.040 370.100 1027.640 432.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.040 1167.600 97.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.040 1167.600 127.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 156.040 1167.600 157.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 186.040 1167.600 187.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 216.040 1167.600 217.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.040 1167.600 247.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 276.040 1167.600 277.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 306.040 1167.600 307.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 336.040 1167.600 337.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 366.040 1167.600 367.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.040 1167.600 397.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 426.040 1167.600 427.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 456.040 1167.600 457.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 486.040 1167.600 487.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 516.040 1167.600 517.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.040 1167.600 547.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 576.040 1167.600 577.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 606.040 1167.600 607.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.040 1167.600 637.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 666.040 1167.600 667.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.040 1167.600 697.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 726.040 1167.600 727.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 756.040 1167.600 757.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.040 1167.600 787.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.040 1167.600 817.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.040 1167.600 847.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 876.040 1167.600 877.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 906.040 1167.600 907.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 936.040 1167.600 937.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 966.040 1167.600 967.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.040 1167.600 997.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1026.040 1167.600 1027.640 1229.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.040 10.640 37.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.040 10.640 67.640 1588.720 ;
    END
  END vssd1
  PIN write_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END write_data[0]
  PIN write_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END write_data[10]
  PIN write_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END write_data[11]
  PIN write_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END write_data[12]
  PIN write_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END write_data[13]
  PIN write_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END write_data[14]
  PIN write_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END write_data[15]
  PIN write_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.080 4.000 376.680 ;
    END
  END write_data[16]
  PIN write_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END write_data[17]
  PIN write_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 4.000 399.800 ;
    END
  END write_data[18]
  PIN write_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END write_data[19]
  PIN write_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END write_data[1]
  PIN write_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 422.320 4.000 422.920 ;
    END
  END write_data[20]
  PIN write_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END write_data[21]
  PIN write_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END write_data[22]
  PIN write_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END write_data[23]
  PIN write_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END write_data[24]
  PIN write_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END write_data[25]
  PIN write_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.680 4.000 492.280 ;
    END
  END write_data[26]
  PIN write_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END write_data[27]
  PIN write_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END write_data[28]
  PIN write_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END write_data[29]
  PIN write_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END write_data[2]
  PIN write_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END write_data[30]
  PIN write_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.160 4.000 550.760 ;
    END
  END write_data[31]
  PIN write_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END write_data[32]
  PIN write_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.280 4.000 573.880 ;
    END
  END write_data[33]
  PIN write_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END write_data[34]
  PIN write_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 596.400 4.000 597.000 ;
    END
  END write_data[35]
  PIN write_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END write_data[36]
  PIN write_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 619.520 4.000 620.120 ;
    END
  END write_data[37]
  PIN write_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END write_data[3]
  PIN write_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END write_data[4]
  PIN write_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END write_data[5]
  PIN write_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END write_data[6]
  PIN write_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END write_data[7]
  PIN write_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END write_data[8]
  PIN write_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END write_data[9]
  PIN write_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END write_en
  OBS
      LAYER li1 ;
        RECT 5.520 1174.275 1050.000 1588.565 ;
        RECT 5.520 379.185 1050.035 1174.275 ;
        RECT 5.520 10.795 1050.000 379.185 ;
      LAYER met1 ;
        RECT 5.520 1149.440 1050.000 1594.380 ;
        RECT 5.520 1147.260 1050.020 1149.440 ;
        RECT 5.520 5.620 1050.000 1147.260 ;
      LAYER met2 ;
        RECT 6.990 1193.770 1050.000 1594.380 ;
        RECT 6.990 275.930 1050.020 1193.770 ;
        RECT 6.990 5.595 1050.000 275.930 ;
      LAYER met3 ;
        RECT 4.000 1060.480 1049.655 1595.000 ;
        RECT 4.400 1059.080 1049.655 1060.480 ;
        RECT 4.000 1048.920 1049.655 1059.080 ;
        RECT 4.400 1047.520 1049.655 1048.920 ;
        RECT 4.000 1037.360 1049.655 1047.520 ;
        RECT 4.400 1035.960 1049.655 1037.360 ;
        RECT 4.000 1025.800 1049.655 1035.960 ;
        RECT 4.400 1024.400 1049.655 1025.800 ;
        RECT 4.000 1014.240 1049.655 1024.400 ;
        RECT 4.400 1012.840 1049.655 1014.240 ;
        RECT 4.000 1002.680 1049.655 1012.840 ;
        RECT 4.400 1001.280 1049.655 1002.680 ;
        RECT 4.000 991.120 1049.655 1001.280 ;
        RECT 4.400 989.720 1049.655 991.120 ;
        RECT 4.000 979.560 1049.655 989.720 ;
        RECT 4.400 978.160 1049.655 979.560 ;
        RECT 4.000 968.000 1049.655 978.160 ;
        RECT 4.400 966.600 1049.655 968.000 ;
        RECT 4.000 956.440 1049.655 966.600 ;
        RECT 4.400 955.040 1049.655 956.440 ;
        RECT 4.000 944.880 1049.655 955.040 ;
        RECT 4.400 943.480 1049.655 944.880 ;
        RECT 4.000 933.320 1049.655 943.480 ;
        RECT 4.400 931.920 1049.655 933.320 ;
        RECT 4.000 921.760 1049.655 931.920 ;
        RECT 4.400 920.360 1049.655 921.760 ;
        RECT 4.000 910.200 1049.655 920.360 ;
        RECT 4.400 908.800 1049.655 910.200 ;
        RECT 4.000 898.640 1049.655 908.800 ;
        RECT 4.400 897.240 1049.655 898.640 ;
        RECT 4.000 887.080 1049.655 897.240 ;
        RECT 4.400 885.680 1049.655 887.080 ;
        RECT 4.000 875.520 1049.655 885.680 ;
        RECT 4.400 874.120 1049.655 875.520 ;
        RECT 4.000 863.960 1049.655 874.120 ;
        RECT 4.400 862.560 1049.655 863.960 ;
        RECT 4.000 852.400 1049.655 862.560 ;
        RECT 4.400 851.000 1049.655 852.400 ;
        RECT 4.000 840.840 1049.655 851.000 ;
        RECT 4.400 839.440 1049.655 840.840 ;
        RECT 4.000 829.280 1049.655 839.440 ;
        RECT 4.400 827.880 1049.655 829.280 ;
        RECT 4.000 817.720 1049.655 827.880 ;
        RECT 4.400 816.320 1049.655 817.720 ;
        RECT 4.000 806.160 1049.655 816.320 ;
        RECT 4.400 804.760 1049.655 806.160 ;
        RECT 4.000 793.920 1049.655 804.760 ;
        RECT 4.400 792.520 1049.655 793.920 ;
        RECT 4.000 782.360 1049.655 792.520 ;
        RECT 4.400 780.960 1049.655 782.360 ;
        RECT 4.000 770.800 1049.655 780.960 ;
        RECT 4.400 769.400 1049.655 770.800 ;
        RECT 4.000 759.240 1049.655 769.400 ;
        RECT 4.400 757.840 1049.655 759.240 ;
        RECT 4.000 747.680 1049.655 757.840 ;
        RECT 4.400 746.280 1049.655 747.680 ;
        RECT 4.000 736.120 1049.655 746.280 ;
        RECT 4.400 734.720 1049.655 736.120 ;
        RECT 4.000 724.560 1049.655 734.720 ;
        RECT 4.400 723.160 1049.655 724.560 ;
        RECT 4.000 713.000 1049.655 723.160 ;
        RECT 4.400 711.600 1049.655 713.000 ;
        RECT 4.000 701.440 1049.655 711.600 ;
        RECT 4.400 700.040 1049.655 701.440 ;
        RECT 4.000 689.880 1049.655 700.040 ;
        RECT 4.400 688.480 1049.655 689.880 ;
        RECT 4.000 678.320 1049.655 688.480 ;
        RECT 4.400 676.920 1049.655 678.320 ;
        RECT 4.000 666.760 1049.655 676.920 ;
        RECT 4.400 665.360 1049.655 666.760 ;
        RECT 4.000 655.200 1049.655 665.360 ;
        RECT 4.400 653.800 1049.655 655.200 ;
        RECT 4.000 643.640 1049.655 653.800 ;
        RECT 4.400 642.240 1049.655 643.640 ;
        RECT 4.000 632.080 1049.655 642.240 ;
        RECT 4.400 630.680 1049.655 632.080 ;
        RECT 4.000 620.520 1049.655 630.680 ;
        RECT 4.400 619.120 1049.655 620.520 ;
        RECT 4.000 608.960 1049.655 619.120 ;
        RECT 4.400 607.560 1049.655 608.960 ;
        RECT 4.000 597.400 1049.655 607.560 ;
        RECT 4.400 596.000 1049.655 597.400 ;
        RECT 4.000 585.840 1049.655 596.000 ;
        RECT 4.400 584.440 1049.655 585.840 ;
        RECT 4.000 574.280 1049.655 584.440 ;
        RECT 4.400 572.880 1049.655 574.280 ;
        RECT 4.000 562.720 1049.655 572.880 ;
        RECT 4.400 561.320 1049.655 562.720 ;
        RECT 4.000 551.160 1049.655 561.320 ;
        RECT 4.400 549.760 1049.655 551.160 ;
        RECT 4.000 539.600 1049.655 549.760 ;
        RECT 4.400 538.200 1049.655 539.600 ;
        RECT 4.000 527.360 1049.655 538.200 ;
        RECT 4.400 525.960 1049.655 527.360 ;
        RECT 4.000 515.800 1049.655 525.960 ;
        RECT 4.400 514.400 1049.655 515.800 ;
        RECT 4.000 504.240 1049.655 514.400 ;
        RECT 4.400 502.840 1049.655 504.240 ;
        RECT 4.000 492.680 1049.655 502.840 ;
        RECT 4.400 491.280 1049.655 492.680 ;
        RECT 4.000 481.120 1049.655 491.280 ;
        RECT 4.400 479.720 1049.655 481.120 ;
        RECT 4.000 469.560 1049.655 479.720 ;
        RECT 4.400 468.160 1049.655 469.560 ;
        RECT 4.000 458.000 1049.655 468.160 ;
        RECT 4.400 456.600 1049.655 458.000 ;
        RECT 4.000 446.440 1049.655 456.600 ;
        RECT 4.400 445.040 1049.655 446.440 ;
        RECT 4.000 434.880 1049.655 445.040 ;
        RECT 4.400 433.480 1049.655 434.880 ;
        RECT 4.000 423.320 1049.655 433.480 ;
        RECT 4.400 421.920 1049.655 423.320 ;
        RECT 4.000 411.760 1049.655 421.920 ;
        RECT 4.400 410.360 1049.655 411.760 ;
        RECT 4.000 400.200 1049.655 410.360 ;
        RECT 4.400 398.800 1049.655 400.200 ;
        RECT 4.000 388.640 1049.655 398.800 ;
        RECT 4.400 387.240 1049.655 388.640 ;
        RECT 4.000 377.080 1049.655 387.240 ;
        RECT 4.400 375.680 1049.655 377.080 ;
        RECT 4.000 365.520 1049.655 375.680 ;
        RECT 4.400 364.120 1049.655 365.520 ;
        RECT 4.000 353.960 1049.655 364.120 ;
        RECT 4.400 352.560 1049.655 353.960 ;
        RECT 4.000 342.400 1049.655 352.560 ;
        RECT 4.400 341.000 1049.655 342.400 ;
        RECT 4.000 330.840 1049.655 341.000 ;
        RECT 4.400 329.440 1049.655 330.840 ;
        RECT 4.000 319.280 1049.655 329.440 ;
        RECT 4.400 317.880 1049.655 319.280 ;
        RECT 4.000 307.720 1049.655 317.880 ;
        RECT 4.400 306.320 1049.655 307.720 ;
        RECT 4.000 296.160 1049.655 306.320 ;
        RECT 4.400 294.760 1049.655 296.160 ;
        RECT 4.000 284.600 1049.655 294.760 ;
        RECT 4.400 283.200 1049.655 284.600 ;
        RECT 4.000 273.040 1049.655 283.200 ;
        RECT 4.400 271.640 1049.655 273.040 ;
        RECT 4.000 260.800 1049.655 271.640 ;
        RECT 4.400 259.400 1049.655 260.800 ;
        RECT 4.000 249.240 1049.655 259.400 ;
        RECT 4.400 247.840 1049.655 249.240 ;
        RECT 4.000 237.680 1049.655 247.840 ;
        RECT 4.400 236.280 1049.655 237.680 ;
        RECT 4.000 226.120 1049.655 236.280 ;
        RECT 4.400 224.720 1049.655 226.120 ;
        RECT 4.000 214.560 1049.655 224.720 ;
        RECT 4.400 213.160 1049.655 214.560 ;
        RECT 4.000 203.000 1049.655 213.160 ;
        RECT 4.400 201.600 1049.655 203.000 ;
        RECT 4.000 191.440 1049.655 201.600 ;
        RECT 4.400 190.040 1049.655 191.440 ;
        RECT 4.000 179.880 1049.655 190.040 ;
        RECT 4.400 178.480 1049.655 179.880 ;
        RECT 4.000 168.320 1049.655 178.480 ;
        RECT 4.400 166.920 1049.655 168.320 ;
        RECT 4.000 156.760 1049.655 166.920 ;
        RECT 4.400 155.360 1049.655 156.760 ;
        RECT 4.000 145.200 1049.655 155.360 ;
        RECT 4.400 143.800 1049.655 145.200 ;
        RECT 4.000 133.640 1049.655 143.800 ;
        RECT 4.400 132.240 1049.655 133.640 ;
        RECT 4.000 122.080 1049.655 132.240 ;
        RECT 4.400 120.680 1049.655 122.080 ;
        RECT 4.000 110.520 1049.655 120.680 ;
        RECT 4.400 109.120 1049.655 110.520 ;
        RECT 4.000 98.960 1049.655 109.120 ;
        RECT 4.400 97.560 1049.655 98.960 ;
        RECT 4.000 87.400 1049.655 97.560 ;
        RECT 4.400 86.000 1049.655 87.400 ;
        RECT 4.000 75.840 1049.655 86.000 ;
        RECT 4.400 74.440 1049.655 75.840 ;
        RECT 4.000 64.280 1049.655 74.440 ;
        RECT 4.400 62.880 1049.655 64.280 ;
        RECT 4.000 52.720 1049.655 62.880 ;
        RECT 4.400 51.320 1049.655 52.720 ;
        RECT 4.000 41.160 1049.655 51.320 ;
        RECT 4.400 39.760 1049.655 41.160 ;
        RECT 4.000 29.600 1049.655 39.760 ;
        RECT 4.400 28.200 1049.655 29.600 ;
        RECT 4.000 18.040 1049.655 28.200 ;
        RECT 4.400 16.640 1049.655 18.040 ;
        RECT 4.000 6.480 1049.655 16.640 ;
        RECT 4.400 5.080 1049.655 6.480 ;
        RECT 4.000 5.000 1049.655 5.080 ;
      LAYER met4 ;
        RECT 11.830 1589.120 1047.090 1595.000 ;
        RECT 11.830 10.240 20.640 1589.120 ;
        RECT 23.040 10.240 35.640 1589.120 ;
        RECT 38.040 10.240 50.640 1589.120 ;
        RECT 53.040 10.240 65.640 1589.120 ;
        RECT 68.040 10.240 80.640 1589.120 ;
        RECT 83.040 1230.300 1047.090 1589.120 ;
        RECT 83.040 1167.200 95.640 1230.300 ;
        RECT 98.040 1167.200 110.640 1230.300 ;
        RECT 113.040 1167.200 125.640 1230.300 ;
        RECT 128.040 1167.200 140.640 1230.300 ;
        RECT 143.040 1167.200 155.640 1230.300 ;
        RECT 158.040 1167.200 170.640 1230.300 ;
        RECT 173.040 1167.200 185.640 1230.300 ;
        RECT 188.040 1167.200 200.640 1230.300 ;
        RECT 203.040 1167.200 215.640 1230.300 ;
        RECT 218.040 1167.200 230.640 1230.300 ;
        RECT 233.040 1167.200 245.640 1230.300 ;
        RECT 248.040 1167.200 260.640 1230.300 ;
        RECT 263.040 1167.200 275.640 1230.300 ;
        RECT 278.040 1167.200 290.640 1230.300 ;
        RECT 293.040 1167.200 305.640 1230.300 ;
        RECT 308.040 1167.200 320.640 1230.300 ;
        RECT 323.040 1167.200 335.640 1230.300 ;
        RECT 338.040 1167.200 350.640 1230.300 ;
        RECT 353.040 1167.200 365.640 1230.300 ;
        RECT 368.040 1167.200 380.640 1230.300 ;
        RECT 383.040 1167.200 395.640 1230.300 ;
        RECT 398.040 1167.200 410.640 1230.300 ;
        RECT 413.040 1167.200 425.640 1230.300 ;
        RECT 428.040 1167.200 440.640 1230.300 ;
        RECT 443.040 1167.200 455.640 1230.300 ;
        RECT 458.040 1167.200 470.640 1230.300 ;
        RECT 473.040 1167.200 485.640 1230.300 ;
        RECT 488.040 1167.200 500.640 1230.300 ;
        RECT 503.040 1167.200 515.640 1230.300 ;
        RECT 518.040 1167.200 530.640 1230.300 ;
        RECT 533.040 1167.200 545.640 1230.300 ;
        RECT 548.040 1167.200 560.640 1230.300 ;
        RECT 563.040 1167.200 575.640 1230.300 ;
        RECT 578.040 1167.200 590.640 1230.300 ;
        RECT 593.040 1167.200 605.640 1230.300 ;
        RECT 608.040 1167.200 620.640 1230.300 ;
        RECT 623.040 1167.200 635.640 1230.300 ;
        RECT 638.040 1167.200 650.640 1230.300 ;
        RECT 653.040 1167.200 665.640 1230.300 ;
        RECT 668.040 1167.200 680.640 1230.300 ;
        RECT 683.040 1167.200 695.640 1230.300 ;
        RECT 698.040 1167.200 710.640 1230.300 ;
        RECT 713.040 1167.200 725.640 1230.300 ;
        RECT 728.040 1167.200 740.640 1230.300 ;
        RECT 743.040 1167.200 755.640 1230.300 ;
        RECT 758.040 1167.200 770.640 1230.300 ;
        RECT 773.040 1167.200 785.640 1230.300 ;
        RECT 788.040 1167.200 800.640 1230.300 ;
        RECT 803.040 1167.200 815.640 1230.300 ;
        RECT 818.040 1167.200 830.640 1230.300 ;
        RECT 833.040 1167.200 845.640 1230.300 ;
        RECT 848.040 1167.200 860.640 1230.300 ;
        RECT 863.040 1167.200 875.640 1230.300 ;
        RECT 878.040 1167.200 890.640 1230.300 ;
        RECT 893.040 1167.200 905.640 1230.300 ;
        RECT 908.040 1167.200 920.640 1230.300 ;
        RECT 923.040 1167.200 935.640 1230.300 ;
        RECT 938.040 1167.200 950.640 1230.300 ;
        RECT 953.040 1167.200 965.640 1230.300 ;
        RECT 968.040 1167.200 980.640 1230.300 ;
        RECT 983.040 1167.200 995.640 1230.300 ;
        RECT 998.040 1167.200 1010.640 1230.300 ;
        RECT 1013.040 1167.200 1025.640 1230.300 ;
        RECT 1028.040 1167.200 1040.640 1230.300 ;
        RECT 1043.040 1167.200 1047.090 1230.300 ;
        RECT 83.040 432.800 1047.090 1167.200 ;
        RECT 83.040 369.700 95.640 432.800 ;
        RECT 98.040 369.700 110.640 432.800 ;
        RECT 113.040 369.700 125.640 432.800 ;
        RECT 128.040 369.700 140.640 432.800 ;
        RECT 143.040 369.700 155.640 432.800 ;
        RECT 158.040 369.700 170.640 432.800 ;
        RECT 173.040 369.700 185.640 432.800 ;
        RECT 188.040 369.700 200.640 432.800 ;
        RECT 203.040 369.700 215.640 432.800 ;
        RECT 218.040 369.700 230.640 432.800 ;
        RECT 233.040 369.700 245.640 432.800 ;
        RECT 248.040 369.700 260.640 432.800 ;
        RECT 263.040 369.700 275.640 432.800 ;
        RECT 278.040 369.700 290.640 432.800 ;
        RECT 293.040 369.700 305.640 432.800 ;
        RECT 308.040 369.700 320.640 432.800 ;
        RECT 323.040 369.700 335.640 432.800 ;
        RECT 338.040 369.700 350.640 432.800 ;
        RECT 353.040 369.700 365.640 432.800 ;
        RECT 368.040 369.700 380.640 432.800 ;
        RECT 383.040 369.700 395.640 432.800 ;
        RECT 398.040 369.700 410.640 432.800 ;
        RECT 413.040 369.700 425.640 432.800 ;
        RECT 428.040 369.700 440.640 432.800 ;
        RECT 443.040 369.700 455.640 432.800 ;
        RECT 458.040 369.700 470.640 432.800 ;
        RECT 473.040 369.700 485.640 432.800 ;
        RECT 488.040 369.700 500.640 432.800 ;
        RECT 503.040 369.700 515.640 432.800 ;
        RECT 518.040 369.700 530.640 432.800 ;
        RECT 533.040 369.700 545.640 432.800 ;
        RECT 548.040 369.700 560.640 432.800 ;
        RECT 563.040 369.700 575.640 432.800 ;
        RECT 578.040 369.700 590.640 432.800 ;
        RECT 593.040 369.700 605.640 432.800 ;
        RECT 608.040 369.700 620.640 432.800 ;
        RECT 623.040 369.700 635.640 432.800 ;
        RECT 638.040 369.700 650.640 432.800 ;
        RECT 653.040 369.700 665.640 432.800 ;
        RECT 668.040 369.700 680.640 432.800 ;
        RECT 683.040 369.700 695.640 432.800 ;
        RECT 698.040 369.700 710.640 432.800 ;
        RECT 713.040 369.700 725.640 432.800 ;
        RECT 728.040 369.700 740.640 432.800 ;
        RECT 743.040 369.700 755.640 432.800 ;
        RECT 758.040 369.700 770.640 432.800 ;
        RECT 773.040 369.700 785.640 432.800 ;
        RECT 788.040 369.700 800.640 432.800 ;
        RECT 803.040 369.700 815.640 432.800 ;
        RECT 818.040 369.700 830.640 432.800 ;
        RECT 833.040 369.700 845.640 432.800 ;
        RECT 848.040 369.700 860.640 432.800 ;
        RECT 863.040 369.700 875.640 432.800 ;
        RECT 878.040 369.700 890.640 432.800 ;
        RECT 893.040 369.700 905.640 432.800 ;
        RECT 908.040 369.700 920.640 432.800 ;
        RECT 923.040 369.700 935.640 432.800 ;
        RECT 938.040 369.700 950.640 432.800 ;
        RECT 953.040 369.700 965.640 432.800 ;
        RECT 968.040 369.700 980.640 432.800 ;
        RECT 983.040 369.700 995.640 432.800 ;
        RECT 998.040 369.700 1010.640 432.800 ;
        RECT 1013.040 369.700 1025.640 432.800 ;
        RECT 1028.040 369.700 1040.640 432.800 ;
        RECT 1043.040 369.700 1047.090 432.800 ;
        RECT 83.040 10.240 1047.090 369.700 ;
        RECT 11.830 5.000 1047.090 10.240 ;
      LAYER met5 ;
        RECT 11.620 439.500 1047.300 1168.700 ;
  END
END sram_38_4096
END LIBRARY

