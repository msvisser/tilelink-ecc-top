VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_32_2048_sky130_mask
   CLASS BLOCK ;
   SIZE 808.9 BY 553.9 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  127.16 0.0 127.54 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  133.96 0.0 134.34 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  138.72 0.0 139.1 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  144.84 0.0 145.22 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  151.64 0.0 152.02 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  156.4 0.0 156.78 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  163.2 0.0 163.58 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  167.96 0.0 168.34 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  174.76 0.0 175.14 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  180.88 0.0 181.26 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  186.32 0.0 186.7 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 0.0 192.82 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  197.88 0.0 198.26 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  204.0 0.0 204.38 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  208.76 0.0 209.14 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  215.56 0.0 215.94 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  221.68 0.0 222.06 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  227.12 0.0 227.5 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  233.24 0.0 233.62 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  238.68 0.0 239.06 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  244.8 0.0 245.18 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  250.92 0.0 251.3 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  256.36 0.0 256.74 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  262.48 0.0 262.86 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  267.24 0.0 267.62 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  274.04 0.0 274.42 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  278.8 0.0 279.18 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  284.92 0.0 285.3 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  291.04 0.0 291.42 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  296.48 0.0 296.86 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  303.28 0.0 303.66 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  308.04 0.0 308.42 1.06 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  314.84 0.0 315.22 1.06 ;
      END
   END din0[32]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  86.36 0.0 86.74 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  92.48 0.0 92.86 1.06 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  97.92 0.0 98.3 1.06 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 175.44 1.06 175.82 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 184.96 1.06 185.34 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 190.4 1.06 190.78 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 199.24 1.06 199.62 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 204.68 1.06 205.06 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 212.84 1.06 213.22 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 218.28 1.06 218.66 ;
      END
   END addr0[9]
   PIN addr0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 227.12 1.06 227.5 ;
      END
   END addr0[10]
   PIN addr0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 231.88 1.06 232.26 ;
      END
   END addr0[11]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 66.64 1.06 67.02 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 75.48 1.06 75.86 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 67.32 1.06 67.7 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.04 0.0 104.42 1.06 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.16 0.0 110.54 1.06 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.28 0.0 116.66 1.06 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  122.4 0.0 122.78 1.06 ;
      END
   END wmask0[3]
   PIN spare_wen0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  320.28 0.0 320.66 1.06 ;
      END
   END spare_wen0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  150.96 0.0 151.34 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.04 0.0 172.42 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  193.12 0.0 193.5 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  212.84 0.0 213.22 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  232.56 0.0 232.94 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  252.96 0.0 253.34 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  271.32 0.0 271.7 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  292.4 0.0 292.78 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  311.44 0.0 311.82 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  332.52 0.0 332.9 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  352.92 0.0 353.3 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  372.64 0.0 373.02 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  393.04 0.0 393.42 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  412.76 0.0 413.14 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  432.48 0.0 432.86 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  452.88 0.0 453.26 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  471.24 0.0 471.62 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  493.0 0.0 493.38 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  512.72 0.0 513.1 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  532.44 0.0 532.82 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  552.84 0.0 553.22 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  572.56 0.0 572.94 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  592.96 0.0 593.34 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  612.68 0.0 613.06 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  633.08 0.0 633.46 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  652.8 0.0 653.18 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  672.52 0.0 672.9 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  692.92 0.0 693.3 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  712.64 0.0 713.02 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  807.84 92.48 808.9 92.86 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  807.84 91.8 808.9 92.18 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  807.84 87.04 808.9 87.42 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  807.84 87.72 808.9 88.1 ;
      END
   END dout0[32]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  4.76 4.76 6.5 550.5 ;
         LAYER met4 ;
         RECT  802.4 4.76 804.14 550.5 ;
         LAYER met3 ;
         RECT  4.76 548.76 804.14 550.5 ;
         LAYER met3 ;
         RECT  4.76 4.76 804.14 6.5 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  805.8 1.36 807.54 553.9 ;
         LAYER met3 ;
         RECT  1.36 552.16 807.54 553.9 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 553.9 ;
         LAYER met3 ;
         RECT  1.36 1.36 807.54 3.1 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 808.28 553.28 ;
   LAYER  met2 ;
      RECT  0.62 0.62 808.28 553.28 ;
   LAYER  met3 ;
      RECT  1.66 174.84 808.28 176.42 ;
      RECT  0.62 176.42 1.66 184.36 ;
      RECT  0.62 185.94 1.66 189.8 ;
      RECT  0.62 191.38 1.66 198.64 ;
      RECT  0.62 200.22 1.66 204.08 ;
      RECT  0.62 205.66 1.66 212.24 ;
      RECT  0.62 213.82 1.66 217.68 ;
      RECT  0.62 219.26 1.66 226.52 ;
      RECT  0.62 228.1 1.66 231.28 ;
      RECT  0.62 76.46 1.66 174.84 ;
      RECT  0.62 68.3 1.66 74.88 ;
      RECT  1.66 91.88 807.24 93.46 ;
      RECT  1.66 93.46 807.24 174.84 ;
      RECT  807.24 93.46 808.28 174.84 ;
      RECT  807.24 88.7 808.28 91.2 ;
      RECT  1.66 176.42 4.16 548.16 ;
      RECT  1.66 548.16 4.16 551.1 ;
      RECT  4.16 176.42 804.74 548.16 ;
      RECT  804.74 176.42 808.28 548.16 ;
      RECT  804.74 548.16 808.28 551.1 ;
      RECT  1.66 4.16 4.16 7.1 ;
      RECT  1.66 7.1 4.16 91.88 ;
      RECT  4.16 7.1 804.74 91.88 ;
      RECT  804.74 4.16 807.24 7.1 ;
      RECT  804.74 7.1 807.24 91.88 ;
      RECT  0.62 232.86 0.76 551.56 ;
      RECT  0.62 551.56 0.76 553.28 ;
      RECT  0.76 232.86 1.66 551.56 ;
      RECT  1.66 551.1 4.16 551.56 ;
      RECT  4.16 551.1 804.74 551.56 ;
      RECT  804.74 551.1 808.14 551.56 ;
      RECT  808.14 551.1 808.28 551.56 ;
      RECT  808.14 551.56 808.28 553.28 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 66.04 ;
      RECT  0.76 0.62 1.66 0.76 ;
      RECT  0.76 3.7 1.66 66.04 ;
      RECT  807.24 0.62 808.14 0.76 ;
      RECT  807.24 3.7 808.14 86.44 ;
      RECT  808.14 0.62 808.28 0.76 ;
      RECT  808.14 0.76 808.28 3.7 ;
      RECT  808.14 3.7 808.28 86.44 ;
      RECT  1.66 0.62 4.16 0.76 ;
      RECT  1.66 3.7 4.16 4.16 ;
      RECT  4.16 0.62 804.74 0.76 ;
      RECT  4.16 3.7 804.74 4.16 ;
      RECT  804.74 0.62 807.24 0.76 ;
      RECT  804.74 3.7 807.24 4.16 ;
   LAYER  met4 ;
      RECT  126.56 1.66 128.14 553.28 ;
      RECT  128.14 0.62 133.36 1.66 ;
      RECT  134.94 0.62 138.12 1.66 ;
      RECT  139.7 0.62 144.24 1.66 ;
      RECT  152.62 0.62 155.8 1.66 ;
      RECT  157.38 0.62 162.6 1.66 ;
      RECT  164.18 0.62 167.36 1.66 ;
      RECT  175.74 0.62 180.28 1.66 ;
      RECT  181.86 0.62 185.72 1.66 ;
      RECT  187.3 0.62 191.84 1.66 ;
      RECT  198.86 0.62 203.4 1.66 ;
      RECT  204.98 0.62 208.16 1.66 ;
      RECT  216.54 0.62 221.08 1.66 ;
      RECT  222.66 0.62 226.52 1.66 ;
      RECT  234.22 0.62 238.08 1.66 ;
      RECT  239.66 0.62 244.2 1.66 ;
      RECT  245.78 0.62 250.32 1.66 ;
      RECT  257.34 0.62 261.88 1.66 ;
      RECT  263.46 0.62 266.64 1.66 ;
      RECT  275.02 0.62 278.2 1.66 ;
      RECT  279.78 0.62 284.32 1.66 ;
      RECT  285.9 0.62 290.44 1.66 ;
      RECT  297.46 0.62 302.68 1.66 ;
      RECT  304.26 0.62 307.44 1.66 ;
      RECT  87.34 0.62 91.88 1.66 ;
      RECT  93.46 0.62 97.32 1.66 ;
      RECT  98.9 0.62 103.44 1.66 ;
      RECT  105.02 0.62 109.56 1.66 ;
      RECT  111.14 0.62 115.68 1.66 ;
      RECT  117.26 0.62 121.8 1.66 ;
      RECT  123.38 0.62 126.56 1.66 ;
      RECT  315.82 0.62 319.68 1.66 ;
      RECT  145.82 0.62 150.36 1.66 ;
      RECT  168.94 0.62 171.44 1.66 ;
      RECT  173.02 0.62 174.16 1.66 ;
      RECT  194.1 0.62 197.28 1.66 ;
      RECT  209.74 0.62 212.24 1.66 ;
      RECT  213.82 0.62 214.96 1.66 ;
      RECT  228.1 0.62 231.96 1.66 ;
      RECT  251.9 0.62 252.36 1.66 ;
      RECT  253.94 0.62 255.76 1.66 ;
      RECT  268.22 0.62 270.72 1.66 ;
      RECT  272.3 0.62 273.44 1.66 ;
      RECT  293.38 0.62 295.88 1.66 ;
      RECT  309.02 0.62 310.84 1.66 ;
      RECT  312.42 0.62 314.24 1.66 ;
      RECT  321.26 0.62 331.92 1.66 ;
      RECT  333.5 0.62 352.32 1.66 ;
      RECT  353.9 0.62 372.04 1.66 ;
      RECT  373.62 0.62 392.44 1.66 ;
      RECT  394.02 0.62 412.16 1.66 ;
      RECT  413.74 0.62 431.88 1.66 ;
      RECT  433.46 0.62 452.28 1.66 ;
      RECT  453.86 0.62 470.64 1.66 ;
      RECT  472.22 0.62 492.4 1.66 ;
      RECT  493.98 0.62 512.12 1.66 ;
      RECT  513.7 0.62 531.84 1.66 ;
      RECT  533.42 0.62 552.24 1.66 ;
      RECT  553.82 0.62 571.96 1.66 ;
      RECT  573.54 0.62 592.36 1.66 ;
      RECT  593.94 0.62 612.08 1.66 ;
      RECT  613.66 0.62 632.48 1.66 ;
      RECT  634.06 0.62 652.2 1.66 ;
      RECT  653.78 0.62 671.92 1.66 ;
      RECT  673.5 0.62 692.32 1.66 ;
      RECT  693.9 0.62 712.04 1.66 ;
      RECT  4.16 1.66 7.1 4.16 ;
      RECT  4.16 551.1 7.1 553.28 ;
      RECT  7.1 1.66 126.56 4.16 ;
      RECT  7.1 4.16 126.56 551.1 ;
      RECT  7.1 551.1 126.56 553.28 ;
      RECT  128.14 1.66 801.8 4.16 ;
      RECT  128.14 4.16 801.8 551.1 ;
      RECT  128.14 551.1 801.8 553.28 ;
      RECT  801.8 1.66 804.74 4.16 ;
      RECT  801.8 551.1 804.74 553.28 ;
      RECT  713.62 0.62 805.2 0.76 ;
      RECT  713.62 0.76 805.2 1.66 ;
      RECT  805.2 0.62 808.14 0.76 ;
      RECT  808.14 0.62 808.28 0.76 ;
      RECT  808.14 0.76 808.28 1.66 ;
      RECT  804.74 1.66 805.2 4.16 ;
      RECT  808.14 1.66 808.28 4.16 ;
      RECT  804.74 4.16 805.2 551.1 ;
      RECT  808.14 4.16 808.28 551.1 ;
      RECT  804.74 551.1 805.2 553.28 ;
      RECT  808.14 551.1 808.28 553.28 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 1.66 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 85.76 0.76 ;
      RECT  3.7 0.76 85.76 1.66 ;
      RECT  0.62 1.66 0.76 4.16 ;
      RECT  3.7 1.66 4.16 4.16 ;
      RECT  0.62 4.16 0.76 551.1 ;
      RECT  3.7 4.16 4.16 551.1 ;
      RECT  0.62 551.1 0.76 553.28 ;
      RECT  3.7 551.1 4.16 553.28 ;
   END
END    sram_32_2048_sky130_mask
END    LIBRARY
