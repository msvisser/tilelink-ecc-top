VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_39_2048_sky130
   CLASS BLOCK ;
   SIZE 959.86 BY 559.34 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.28 0.0 116.66 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  122.4 0.0 122.78 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  127.16 0.0 127.54 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  133.96 0.0 134.34 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  138.72 0.0 139.1 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  145.52 0.0 145.9 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  150.28 0.0 150.66 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  156.4 0.0 156.78 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  163.2 0.0 163.58 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  168.64 0.0 169.02 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  174.08 0.0 174.46 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  180.2 0.0 180.58 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  185.64 0.0 186.02 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 0.0 192.82 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  197.2 0.0 197.58 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  204.0 0.0 204.38 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  208.76 0.0 209.14 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  215.56 0.0 215.94 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  221.68 0.0 222.06 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  227.12 0.0 227.5 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  232.56 0.0 232.94 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  238.68 0.0 239.06 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  244.8 0.0 245.18 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  250.24 0.0 250.62 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  256.36 0.0 256.74 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  262.48 0.0 262.86 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  267.24 0.0 267.62 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  274.04 0.0 274.42 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  278.8 0.0 279.18 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  285.6 0.0 285.98 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  291.04 0.0 291.42 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  297.16 0.0 297.54 1.06 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  302.6 0.0 302.98 1.06 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  308.72 0.0 309.1 1.06 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  314.16 0.0 314.54 1.06 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  320.28 0.0 320.66 1.06 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  325.72 0.0 326.1 1.06 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  332.52 0.0 332.9 1.06 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  337.28 0.0 337.66 1.06 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  344.08 0.0 344.46 1.06 ;
      END
   END din0[39]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  98.6 0.0 98.98 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.72 0.0 105.1 1.06 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.16 0.0 110.54 1.06 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 180.88 1.06 181.26 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 190.4 1.06 190.78 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 196.52 1.06 196.9 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 204.68 1.06 205.06 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 210.12 1.06 210.5 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 218.28 1.06 218.66 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 223.72 1.06 224.1 ;
      END
   END addr0[9]
   PIN addr0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 232.56 1.06 232.94 ;
      END
   END addr0[10]
   PIN addr0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 238.68 1.06 239.06 ;
      END
   END addr0[11]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 72.08 1.06 72.46 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 80.24 1.06 80.62 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 72.76 1.06 73.14 ;
      END
   END clk0
   PIN spare_wen0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  349.52 0.0 349.9 1.06 ;
      END
   END spare_wen0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  163.88 0.0 164.26 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  183.6 0.0 183.98 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.68 0.0 205.06 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  224.4 0.0 224.78 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  244.12 0.0 244.5 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  264.52 0.0 264.9 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  282.88 0.0 283.26 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  303.96 0.0 304.34 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  323.68 0.0 324.06 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  343.4 0.0 343.78 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  364.48 0.0 364.86 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  384.2 0.0 384.58 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  404.6 0.0 404.98 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  424.32 0.0 424.7 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  444.04 0.0 444.42 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  464.44 0.0 464.82 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  484.16 0.0 484.54 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  504.56 0.0 504.94 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  524.28 0.0 524.66 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  544.0 0.0 544.38 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  564.4 0.0 564.78 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  584.12 0.0 584.5 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  604.52 0.0 604.9 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  624.24 0.0 624.62 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  644.64 0.0 645.02 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  664.36 0.0 664.74 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  684.08 0.0 684.46 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  704.48 0.0 704.86 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  724.2 0.0 724.58 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  744.6 0.0 744.98 1.06 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  764.32 0.0 764.7 1.06 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  784.72 0.0 785.1 1.06 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  804.44 0.0 804.82 1.06 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  824.16 0.0 824.54 1.06 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  844.56 0.0 844.94 1.06 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  864.28 0.0 864.66 1.06 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  958.8 97.24 959.86 97.62 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  958.8 92.48 959.86 92.86 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  958.8 93.16 959.86 93.54 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  958.8 93.84 959.86 94.22 ;
      END
   END dout0[39]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  4.76 554.2 955.1 555.94 ;
         LAYER met3 ;
         RECT  4.76 4.76 955.1 6.5 ;
         LAYER met4 ;
         RECT  4.76 4.76 6.5 555.94 ;
         LAYER met4 ;
         RECT  953.36 4.76 955.1 555.94 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  956.76 1.36 958.5 559.34 ;
         LAYER met3 ;
         RECT  1.36 1.36 958.5 3.1 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 559.34 ;
         LAYER met3 ;
         RECT  1.36 557.6 958.5 559.34 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 959.24 558.72 ;
   LAYER  met2 ;
      RECT  0.62 0.62 959.24 558.72 ;
   LAYER  met3 ;
      RECT  1.66 180.28 959.24 181.86 ;
      RECT  0.62 181.86 1.66 189.8 ;
      RECT  0.62 191.38 1.66 195.92 ;
      RECT  0.62 197.5 1.66 204.08 ;
      RECT  0.62 205.66 1.66 209.52 ;
      RECT  0.62 211.1 1.66 217.68 ;
      RECT  0.62 219.26 1.66 223.12 ;
      RECT  0.62 224.7 1.66 231.96 ;
      RECT  0.62 233.54 1.66 238.08 ;
      RECT  0.62 81.22 1.66 180.28 ;
      RECT  0.62 73.74 1.66 79.64 ;
      RECT  1.66 96.64 958.2 98.22 ;
      RECT  1.66 98.22 958.2 180.28 ;
      RECT  958.2 98.22 959.24 180.28 ;
      RECT  958.2 94.82 959.24 96.64 ;
      RECT  1.66 181.86 4.16 553.6 ;
      RECT  1.66 553.6 4.16 556.54 ;
      RECT  4.16 181.86 955.7 553.6 ;
      RECT  955.7 181.86 959.24 553.6 ;
      RECT  955.7 553.6 959.24 556.54 ;
      RECT  1.66 4.16 4.16 7.1 ;
      RECT  1.66 7.1 4.16 96.64 ;
      RECT  4.16 7.1 955.7 96.64 ;
      RECT  955.7 4.16 958.2 7.1 ;
      RECT  955.7 7.1 958.2 96.64 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 71.48 ;
      RECT  0.76 0.62 1.66 0.76 ;
      RECT  0.76 3.7 1.66 71.48 ;
      RECT  958.2 0.62 959.1 0.76 ;
      RECT  958.2 3.7 959.1 91.88 ;
      RECT  959.1 0.62 959.24 0.76 ;
      RECT  959.1 0.76 959.24 3.7 ;
      RECT  959.1 3.7 959.24 91.88 ;
      RECT  1.66 0.62 4.16 0.76 ;
      RECT  1.66 3.7 4.16 4.16 ;
      RECT  4.16 0.62 955.7 0.76 ;
      RECT  4.16 3.7 955.7 4.16 ;
      RECT  955.7 0.62 958.2 0.76 ;
      RECT  955.7 3.7 958.2 4.16 ;
      RECT  0.62 239.66 0.76 557.0 ;
      RECT  0.62 557.0 0.76 558.72 ;
      RECT  0.76 239.66 1.66 557.0 ;
      RECT  1.66 556.54 4.16 557.0 ;
      RECT  4.16 556.54 955.7 557.0 ;
      RECT  955.7 556.54 959.1 557.0 ;
      RECT  959.1 556.54 959.24 557.0 ;
      RECT  959.1 557.0 959.24 558.72 ;
   LAYER  met4 ;
      RECT  115.68 1.66 117.26 558.72 ;
      RECT  117.26 0.62 121.8 1.66 ;
      RECT  123.38 0.62 126.56 1.66 ;
      RECT  128.14 0.62 133.36 1.66 ;
      RECT  134.94 0.62 138.12 1.66 ;
      RECT  139.7 0.62 144.92 1.66 ;
      RECT  146.5 0.62 149.68 1.66 ;
      RECT  151.26 0.62 155.8 1.66 ;
      RECT  157.38 0.62 162.6 1.66 ;
      RECT  169.62 0.62 173.48 1.66 ;
      RECT  175.06 0.62 179.6 1.66 ;
      RECT  186.62 0.62 191.84 1.66 ;
      RECT  193.42 0.62 196.6 1.66 ;
      RECT  198.18 0.62 203.4 1.66 ;
      RECT  209.74 0.62 214.96 1.66 ;
      RECT  216.54 0.62 221.08 1.66 ;
      RECT  228.1 0.62 231.96 1.66 ;
      RECT  233.54 0.62 238.08 1.66 ;
      RECT  245.78 0.62 249.64 1.66 ;
      RECT  251.22 0.62 255.76 1.66 ;
      RECT  257.34 0.62 261.88 1.66 ;
      RECT  268.22 0.62 273.44 1.66 ;
      RECT  275.02 0.62 278.2 1.66 ;
      RECT  286.58 0.62 290.44 1.66 ;
      RECT  292.02 0.62 296.56 1.66 ;
      RECT  298.14 0.62 302.0 1.66 ;
      RECT  309.7 0.62 313.56 1.66 ;
      RECT  315.14 0.62 319.68 1.66 ;
      RECT  326.7 0.62 331.92 1.66 ;
      RECT  333.5 0.62 336.68 1.66 ;
      RECT  99.58 0.62 104.12 1.66 ;
      RECT  105.7 0.62 109.56 1.66 ;
      RECT  111.14 0.62 115.68 1.66 ;
      RECT  345.06 0.62 348.92 1.66 ;
      RECT  164.86 0.62 168.04 1.66 ;
      RECT  181.18 0.62 183.0 1.66 ;
      RECT  184.58 0.62 185.04 1.66 ;
      RECT  205.66 0.62 208.16 1.66 ;
      RECT  222.66 0.62 223.8 1.66 ;
      RECT  225.38 0.62 226.52 1.66 ;
      RECT  239.66 0.62 243.52 1.66 ;
      RECT  263.46 0.62 263.92 1.66 ;
      RECT  265.5 0.62 266.64 1.66 ;
      RECT  279.78 0.62 282.28 1.66 ;
      RECT  283.86 0.62 285.0 1.66 ;
      RECT  304.94 0.62 308.12 1.66 ;
      RECT  321.26 0.62 323.08 1.66 ;
      RECT  324.66 0.62 325.12 1.66 ;
      RECT  338.26 0.62 342.8 1.66 ;
      RECT  350.5 0.62 363.88 1.66 ;
      RECT  365.46 0.62 383.6 1.66 ;
      RECT  385.18 0.62 404.0 1.66 ;
      RECT  405.58 0.62 423.72 1.66 ;
      RECT  425.3 0.62 443.44 1.66 ;
      RECT  445.02 0.62 463.84 1.66 ;
      RECT  465.42 0.62 483.56 1.66 ;
      RECT  485.14 0.62 503.96 1.66 ;
      RECT  505.54 0.62 523.68 1.66 ;
      RECT  525.26 0.62 543.4 1.66 ;
      RECT  544.98 0.62 563.8 1.66 ;
      RECT  565.38 0.62 583.52 1.66 ;
      RECT  585.1 0.62 603.92 1.66 ;
      RECT  605.5 0.62 623.64 1.66 ;
      RECT  625.22 0.62 644.04 1.66 ;
      RECT  645.62 0.62 663.76 1.66 ;
      RECT  665.34 0.62 683.48 1.66 ;
      RECT  685.06 0.62 703.88 1.66 ;
      RECT  705.46 0.62 723.6 1.66 ;
      RECT  725.18 0.62 744.0 1.66 ;
      RECT  745.58 0.62 763.72 1.66 ;
      RECT  765.3 0.62 784.12 1.66 ;
      RECT  785.7 0.62 803.84 1.66 ;
      RECT  805.42 0.62 823.56 1.66 ;
      RECT  825.14 0.62 843.96 1.66 ;
      RECT  845.54 0.62 863.68 1.66 ;
      RECT  4.16 1.66 7.1 4.16 ;
      RECT  4.16 556.54 7.1 558.72 ;
      RECT  7.1 1.66 115.68 4.16 ;
      RECT  7.1 4.16 115.68 556.54 ;
      RECT  7.1 556.54 115.68 558.72 ;
      RECT  117.26 1.66 952.76 4.16 ;
      RECT  117.26 4.16 952.76 556.54 ;
      RECT  117.26 556.54 952.76 558.72 ;
      RECT  952.76 1.66 955.7 4.16 ;
      RECT  952.76 556.54 955.7 558.72 ;
      RECT  865.26 0.62 956.16 0.76 ;
      RECT  865.26 0.76 956.16 1.66 ;
      RECT  956.16 0.62 959.1 0.76 ;
      RECT  959.1 0.62 959.24 0.76 ;
      RECT  959.1 0.76 959.24 1.66 ;
      RECT  955.7 1.66 956.16 4.16 ;
      RECT  959.1 1.66 959.24 4.16 ;
      RECT  955.7 4.16 956.16 556.54 ;
      RECT  959.1 4.16 959.24 556.54 ;
      RECT  955.7 556.54 956.16 558.72 ;
      RECT  959.1 556.54 959.24 558.72 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 1.66 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 98.0 0.76 ;
      RECT  3.7 0.76 98.0 1.66 ;
      RECT  0.62 1.66 0.76 4.16 ;
      RECT  3.7 1.66 4.16 4.16 ;
      RECT  0.62 4.16 0.76 556.54 ;
      RECT  3.7 4.16 4.16 556.54 ;
      RECT  0.62 556.54 0.76 558.72 ;
      RECT  3.7 556.54 4.16 558.72 ;
   END
END    sram_39_2048_sky130
END    LIBRARY
